netcdf o {
dimensions:
	t = UNLIMITED ; // (31 currently)
	x = 20 ;
	y = 20 ;
variables:
	float t(t) ;
		t:long_name = "Time" ;
		t:units = "seconds since simulation start" ;
	float x(x) ;
	float y(y) ;
	float t_max ;
	float l_boundary ;
	float r_boundary ;
	float t_boundary ;
	float b_boundary ;
	float h(t, y, x) ;
	float hu(t, y, x) ;
	float hv(t, y, x) ;
	float b(y, x) ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:title = "Computed tsunami solution" ;
		:history = "SWE" ;
		:institution = "Technische Universitaet Muenchen, Department of Informatics, Chair of Scientific Computing" ;
		:source = "Bathymetry and displacement data." ;
		:references = "http://www5.in.tum.de/SWE" ;
		:comment = "SWE is free software and licensed under the GNU General Public License. Remark: In general this does not hold for the used input data." ;
data:

 t = 0, 0.2287608, 0.3674662, 0.500887, 0.6985019, 0.8988496, 1.035777, 
    1.172752, 1.376863, 1.513404, 1.721124, 1.861454, 2.002371, 2.215259, 
    2.357662, 2.500283, 2.714231, 2.856667, 3.070328, 3.213333, 3.356624, 
    3.500261, 3.717091, 3.862081, 4.007576, 4.227118, 4.374319, 4.521488, 
    4.668321, 4.887586, 5.032344 ;

 x = 2.25, 6.75, 11.25, 15.75, 20.25, 24.75, 29.25, 33.75, 38.25, 42.75, 
    47.25, 51.75, 56.25, 60.75, 65.25, 69.75, 74.25, 78.75, 83.25, 87.75 ;

 y = 2.25, 6.75, 11.25, 15.75, 20.25, 24.75, 29.25, 33.75, 38.25, 42.75, 
    47.25, 51.75, 56.25, 60.75, 65.25, 69.75, 74.25, 78.75, 83.25, 87.75 ;

 t_max = 100 ;

 l_boundary = 1 ;

 r_boundary = 1 ;

 t_boundary = 1 ;

 b_boundary = 1 ;

 h =
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50, 50.00089, 50.01964, 50.14318, 50.39871, 50.54031, 50.56227, 
    50.5633, 50.5633, 50.5633, 50.5633, 50.5633, 50.56227, 50.54031, 
    50.39871, 50.14318, 50.01964, 50.00089,
  50, 50, 50, 50.01914, 50.21582, 50.95889, 52.25088, 53.0721, 53.28872, 
    53.31026, 53.31026, 53.31026, 53.31026, 53.31026, 53.28872, 53.0721, 
    52.25088, 50.95889, 50.21582, 50.01914,
  50, 50, 50, 50.14206, 50.94887, 52.61259, 54.74611, 56.51145, 57.28546, 
    57.41597, 57.41597, 57.41597, 57.41597, 57.41597, 57.28546, 56.51145, 
    54.74611, 52.61259, 50.94887, 50.14206,
  50, 50, 50, 50.41703, 52.33274, 54.80562, 37.16891, 40.10178, 41.85542, 
    42.20115, 42.20115, 42.20115, 42.20115, 42.20115, 41.85542, 40.10178, 
    37.16891, 54.80562, 52.33274, 50.41703,
  50, 50, 50, 50.543, 53.08184, 56.46067, 40.16543, 44.23988, 46.53956, 
    46.99757, 46.99757, 46.99757, 46.99757, 46.99757, 46.53956, 44.23988, 
    40.16543, 56.46067, 53.08184, 50.543,
  50, 50, 50, 50.56236, 53.28883, 57.26506, 41.88169, 46.54629, 49.0268, 
    49.51175, 49.51175, 49.51175, 49.51175, 49.51175, 49.0268, 46.54629, 
    41.88169, 57.26506, 53.28883, 50.56236,
  50, 50, 50, 50.5633, 53.31026, 57.41597, 42.20115, 46.99757, 49.51175, 50, 
    50, 50, 50, 50, 49.51175, 46.99757, 42.20115, 57.41597, 53.31026, 50.5633,
  50, 50, 50, 50.5633, 53.31026, 57.41597, 42.20115, 46.99757, 49.51175, 50, 
    50, 50, 50, 50, 49.51175, 46.99757, 42.20115, 57.41597, 53.31026, 50.5633,
  50, 50, 50, 50.5633, 53.31026, 57.41597, 42.20115, 46.99757, 49.51175, 50, 
    50, 50, 50, 50, 49.51175, 46.99757, 42.20115, 57.41597, 53.31026, 50.5633,
  50, 50, 50, 50.5633, 53.31026, 57.41597, 42.20115, 46.99757, 49.51175, 50, 
    50, 50, 50, 50, 49.51175, 46.99757, 42.20115, 57.41597, 53.31026, 50.5633,
  50, 50, 50, 50.5633, 53.31026, 57.41597, 42.20115, 46.99757, 49.51175, 50, 
    50, 50, 50, 50, 49.51175, 46.99757, 42.20115, 57.41597, 53.31026, 50.5633,
  50, 50, 50, 50.56236, 53.28883, 57.26506, 41.88169, 46.54629, 49.0268, 
    49.51175, 49.51175, 49.51175, 49.51175, 49.51175, 49.0268, 46.54629, 
    41.88169, 57.26506, 53.28883, 50.56236,
  50, 50, 50, 50.543, 53.08184, 56.46067, 40.16543, 44.23988, 46.53956, 
    46.99757, 46.99757, 46.99757, 46.99757, 46.99757, 46.53956, 44.23988, 
    40.16543, 56.46067, 53.08184, 50.543,
  50, 50, 50, 50.41703, 52.33274, 54.80562, 37.16891, 40.10178, 41.85542, 
    42.20115, 42.20115, 42.20115, 42.20115, 42.20115, 41.85542, 40.10178, 
    37.16891, 54.80562, 52.33274, 50.41703,
  50, 50, 50, 50.14206, 50.94887, 52.61259, 54.74611, 56.51145, 57.28546, 
    57.41597, 57.41597, 57.41597, 57.41597, 57.41597, 57.28546, 56.51145, 
    54.74611, 52.61259, 50.94887, 50.14206,
  50, 50, 50, 50.01914, 50.21582, 50.95889, 52.25088, 53.0721, 53.28872, 
    53.31026, 53.31026, 53.31026, 53.31026, 53.31026, 53.28872, 53.0721, 
    52.25088, 50.95889, 50.21582, 50.01914,
  50, 50, 50, 50.00089, 50.01964, 50.14318, 50.39871, 50.54031, 50.56227, 
    50.5633, 50.5633, 50.5633, 50.5633, 50.5633, 50.56227, 50.54031, 
    50.39871, 50.14318, 50.01964, 50.00089,
  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
  50, 50, 50.00003, 50.00052, 50.00433, 50.01921, 50.04509, 50.06191, 
    50.06643, 50.06701, 50.06704, 50.06705, 50.06704, 50.06701, 50.06643, 
    50.06191, 50.04509, 50.01921, 50.00433, 50.00055,
  50, 50.00003, 50.00087, 50.00961, 50.05626, 50.20186, 50.44462, 50.61497, 
    50.67217, 50.68303, 50.68407, 50.6841, 50.68407, 50.68303, 50.67217, 
    50.61497, 50.44462, 50.20186, 50.0563, 50.01047,
  50, 50.0005, 50.00954, 50.07364, 50.31868, 50.90077, 51.77998, 52.45498, 
    52.74399, 52.81998, 52.83086, 52.83147, 52.83086, 52.81998, 52.74399, 
    52.45498, 51.77998, 50.90077, 50.31919, 50.08321,
  50, 50.00425, 50.0561, 50.31994, 51.04209, 52.23935, 53.72222, 55.04995, 
    55.80231, 56.06958, 56.12353, 56.12822, 56.12353, 56.06958, 55.80231, 
    55.04995, 53.72222, 52.23935, 51.04639, 50.37642,
  50, 50.01937, 50.2041, 50.90802, 52.23825, 53.59549, 54.77774, 56.38982, 
    57.67819, 58.28198, 58.43776, 58.45448, 58.43776, 58.28198, 57.67819, 
    56.38982, 54.77774, 53.59549, 52.2578, 51.1137,
  50, 50.04689, 50.46362, 51.85099, 53.82918, 54.85673, 34.85571, 36.76944, 
    38.87077, 39.97232, 40.2774, 40.31147, 40.2774, 39.97232, 38.87077, 
    36.76944, 34.85571, 54.85673, 53.87556, 52.31464,
  50, 50.06253, 50.62127, 52.47569, 55.05963, 56.32131, 36.81181, 39.63404, 
    42.4338, 43.88548, 44.29691, 44.34454, 44.29691, 43.88548, 42.4338, 
    39.63404, 36.81181, 56.32131, 55.12132, 53.09667,
  50, 50.0665, 50.67325, 52.7473, 55.79268, 57.60468, 38.9283, 42.45947, 
    45.64072, 47.25572, 47.71408, 47.76778, 47.71408, 47.25572, 45.64072, 
    42.45947, 38.9283, 57.60468, 55.85838, 53.42085,
  50, 50.06701, 50.68312, 52.82023, 56.0658, 58.25498, 39.99784, 43.8993, 
    47.2587, 48.93759, 49.41123, 49.46668, 49.41123, 48.93759, 47.2587, 
    43.8993, 39.99784, 58.25499, 56.13206, 53.504,
  50, 50.06705, 50.68407, 52.83086, 56.12307, 58.434, 40.28124, 44.2992, 
    47.71473, 49.41132, 49.88843, 49.9442, 49.88843, 49.41132, 47.71473, 
    44.2992, 40.28124, 58.43401, 56.18938, 53.51565,
  50, 50.06705, 50.6841, 52.83147, 56.12822, 58.45448, 40.31147, 44.34454, 
    47.76778, 49.46668, 49.9442, 50, 49.9442, 49.46668, 47.76778, 44.34454, 
    40.31147, 58.45448, 56.19454, 53.5163,
  50, 50.06705, 50.68407, 52.83086, 56.12307, 58.434, 40.28124, 44.2992, 
    47.71473, 49.41132, 49.88843, 49.9442, 49.88843, 49.41132, 47.71473, 
    44.2992, 40.28124, 58.43401, 56.18938, 53.51565,
  50, 50.06701, 50.68312, 52.82023, 56.0658, 58.25498, 39.99784, 43.8993, 
    47.2587, 48.93759, 49.41123, 49.46668, 49.41123, 48.93759, 47.2587, 
    43.8993, 39.99784, 58.25499, 56.13206, 53.504,
  50, 50.0665, 50.67325, 52.7473, 55.79268, 57.60468, 38.9283, 42.45947, 
    45.64072, 47.25572, 47.71408, 47.76778, 47.71408, 47.25572, 45.64072, 
    42.45947, 38.9283, 57.60468, 55.85838, 53.42085,
  50, 50.06253, 50.62127, 52.47569, 55.05963, 56.32131, 36.81181, 39.63404, 
    42.4338, 43.88548, 44.29691, 44.34454, 44.29691, 43.88548, 42.4338, 
    39.63404, 36.81181, 56.32131, 55.12132, 53.09667,
  50, 50.04689, 50.46362, 51.85099, 53.82918, 54.85673, 34.85571, 36.76944, 
    38.87077, 39.97232, 40.2774, 40.31147, 40.2774, 39.97232, 38.87077, 
    36.76944, 34.85571, 54.85673, 53.87556, 52.31464,
  50, 50.01937, 50.2041, 50.90802, 52.23825, 53.59549, 54.77774, 56.38982, 
    57.67819, 58.28198, 58.43776, 58.45448, 58.43776, 58.28198, 57.67819, 
    56.38982, 54.77774, 53.59549, 52.2578, 51.1137,
  50, 50.00425, 50.05611, 50.32022, 51.04542, 52.25745, 53.76792, 55.1123, 
    55.86828, 56.13589, 56.18985, 56.19454, 56.18985, 56.13589, 55.86828, 
    55.1123, 53.76792, 52.25745, 51.04972, 50.3767,
  50, 50.0005, 50.00981, 50.07932, 50.3634, 51.09147, 52.23401, 53.08366, 
    53.42159, 53.50447, 53.51569, 53.5163, 53.51569, 53.50447, 53.42159, 
    53.08366, 52.23401, 51.09147, 50.36391, 50.08916,
  50, 50.00003, 50.00035, 50.00248, 50.01135, 50.03508, 50.07144, 50.09849, 
    50.10925, 50.11189, 50.1123, 50.11233, 50.1123, 50.11189, 50.10925, 
    50.09849, 50.07144, 50.03508, 50.01138, 50.00283,
  50.00003, 50.00047, 50.00397, 50.02144, 50.07945, 50.21272, 50.41058, 
    50.56773, 50.64073, 50.6633, 50.66787, 50.6684, 50.66787, 50.6633, 
    50.64073, 50.56773, 50.41058, 50.21275, 50.07992, 50.02542,
  50.00035, 50.00396, 50.02623, 50.1137, 50.34717, 50.79665, 51.42458, 
    51.957, 52.2456, 52.35545, 52.38384, 52.38808, 52.38384, 52.35545, 
    52.2456, 51.957, 51.4246, 50.797, 50.3512, 50.14013,
  50.00248, 50.02142, 50.11395, 50.40117, 51.00323, 51.91445, 53.04183, 
    54.08997, 54.76888, 55.08762, 55.19177, 55.21125, 55.19177, 55.08762, 
    54.76888, 54.08997, 53.04195, 51.9169, 51.02522, 50.51666,
  50.01144, 50.07999, 50.35038, 51.00994, 52.04915, 53.17754, 54.30956, 
    55.61894, 56.68689, 57.3087, 57.56064, 57.61737, 57.56064, 57.3087, 
    56.68689, 55.61894, 54.31022, 53.18854, 52.131, 51.36608,
  50.03579, 50.21677, 50.80981, 51.93235, 53.18, 54.02256, 54.54498, 
    55.76036, 57.1125, 58.08554, 58.55375, 58.67302, 58.55375, 58.08554, 
    57.1125, 55.76036, 54.54707, 54.05557, 53.39859, 52.75272,
  50.07394, 50.42658, 51.4799, 53.14213, 54.41399, 54.64256, 33.83235, 
    34.89952, 36.73234, 38.20626, 38.95488, 39.1509, 38.95488, 38.20626, 
    36.73234, 34.89952, 33.83651, 54.70812, 54.83619, 54.62944,
  50.09967, 50.57544, 51.98136, 54.12177, 55.61962, 55.71009, 34.91116, 
    36.62406, 39.12669, 41.05417, 42.03593, 42.29757, 42.03593, 41.05417, 
    39.12669, 36.62406, 34.91661, 55.79733, 56.18638, 56.11113,
  50.10953, 50.64294, 52.2526, 54.77235, 56.65668, 57.01479, 36.78143, 
    39.15889, 42.10759, 44.29716, 45.41027, 45.70964, 45.41027, 44.29716, 
    42.10759, 39.15889, 36.78729, 57.11048, 57.28955, 57.03507,
  50.11193, 50.6637, 52.3568, 55.08623, 57.28836, 58.01969, 38.25213, 
    41.08711, 44.30775, 46.64122, 47.81941, 48.13638, 47.81941, 46.64122, 
    44.30775, 41.08711, 38.25811, 58.11765, 57.94254, 57.4566,
  50.1123, 50.66792, 52.384, 55.19103, 57.5533, 58.52791, 38.97588, 42.05181, 
    45.41687, 47.82088, 49.027, 49.35072, 49.027, 47.82088, 45.41687, 
    42.05181, 38.98189, 58.62634, 58.21232, 57.59066,
  50.11233, 50.66841, 52.3881, 55.21097, 57.61458, 58.66226, 39.16013, 
    42.30486, 45.71302, 48.13736, 49.35086, 49.67621, 49.35086, 48.13736, 
    45.71302, 42.30486, 39.16614, 58.76077, 58.2743, 57.61522,
  50.1123, 50.66792, 52.384, 55.19103, 57.5533, 58.52791, 38.97588, 42.05181, 
    45.41687, 47.82088, 49.027, 49.35072, 49.027, 47.82088, 45.41687, 
    42.05181, 38.98189, 58.62634, 58.21232, 57.59066,
  50.11193, 50.6637, 52.3568, 55.08623, 57.28836, 58.01969, 38.25213, 
    41.08711, 44.30775, 46.64122, 47.81941, 48.13638, 47.81941, 46.64122, 
    44.30775, 41.08711, 38.25811, 58.11765, 57.94254, 57.4566,
  50.10953, 50.64294, 52.2526, 54.77235, 56.65668, 57.01479, 36.78143, 
    39.15889, 42.10759, 44.29716, 45.41027, 45.70964, 45.41027, 44.29716, 
    42.10759, 39.15889, 36.78729, 57.11048, 57.28955, 57.03507,
  50.09967, 50.57544, 51.98136, 54.12177, 55.61962, 55.71009, 34.91116, 
    36.62406, 39.12669, 41.05416, 42.03593, 42.29757, 42.03593, 41.05416, 
    39.12669, 36.62406, 34.91661, 55.79733, 56.18638, 56.11113,
  50.07394, 50.42658, 51.47991, 53.14221, 54.41455, 54.64465, 33.83652, 
    34.90501, 36.73824, 38.21225, 38.96089, 39.15691, 38.96089, 38.21225, 
    36.73824, 34.90501, 33.84068, 54.71021, 54.83675, 54.62954,
  50.03579, 50.21678, 50.81002, 51.93414, 53.18938, 54.05386, 54.60996, 
    55.84837, 57.20882, 58.18375, 58.65225, 58.77155, 58.65225, 58.18375, 
    57.20882, 55.84837, 54.61205, 54.08687, 53.40799, 52.75472,
  50.01144, 50.08019, 50.35281, 51.0263, 52.1191, 53.38277, 54.7231, 
    56.19058, 57.32518, 57.96517, 58.22022, 58.27725, 58.22022, 57.96517, 
    57.32518, 56.19058, 54.72376, 53.39378, 52.20115, 51.38488,
  50.00256, 50.02317, 50.13047, 50.48958, 51.31209, 52.68647, 54.49187, 
    56.10179, 57.0595, 57.47086, 57.59464, 57.61635, 57.59464, 57.47086, 
    57.0595, 56.10179, 54.49199, 52.689, 51.33589, 50.62177,
  50.00129, 50.0064, 50.02679, 50.08691, 50.22361, 50.46659, 50.79207, 
    51.08068, 51.25708, 51.338, 51.36597, 51.37192, 51.36597, 51.338, 
    51.25708, 51.08069, 50.79223, 50.46778, 50.23015, 50.11397,
  50.00669, 50.02701, 50.0945, 50.25881, 50.56988, 51.04548, 51.64762, 
    52.21279, 52.60438, 52.81677, 52.90512, 52.927, 52.90512, 52.81677, 
    52.60439, 52.21289, 51.64861, 51.05164, 50.59788, 50.35524,
  50.02785, 50.09489, 50.28588, 50.67601, 51.28914, 52.07408, 52.98506, 
    53.89861, 54.61225, 55.06088, 55.27913, 55.34003, 55.27913, 55.06088, 
    54.61229, 53.89919, 52.98967, 52.09921, 51.38817, 50.97035,
  50.08994, 50.26125, 50.67938, 51.38288, 52.26771, 53.16558, 54.07648, 
    55.13085, 56.09232, 56.79818, 57.19645, 57.31977, 57.19645, 56.79819, 
    56.09252, 55.13314, 54.09261, 53.24335, 52.53808, 52.08428,
  50.23071, 50.57903, 51.30367, 52.28044, 53.21305, 53.90401, 54.4489, 
    55.38418, 56.44826, 57.36977, 57.96286, 58.1623, 57.96286, 57.3698, 
    56.44889, 55.39082, 54.49197, 54.09322, 53.80024, 53.61964,
  50.48051, 51.06798, 52.10405, 53.18523, 53.90469, 54.21851, 54.2399, 
    54.91967, 55.99562, 57.10949, 57.91224, 58.19943, 57.91224, 57.10954, 
    55.99687, 54.93334, 54.32989, 54.59401, 54.96481, 55.33045,
  50.81744, 51.70311, 53.0743, 54.17511, 54.54577, 54.3563, 33.30655, 
    33.55083, 34.69957, 36.12558, 37.21526, 37.61398, 37.21526, 36.12564, 
    34.70108, 33.57091, 33.46097, 54.97598, 56.21574, 57.30429,
  51.09428, 52.24483, 53.93998, 55.15546, 55.38615, 54.91632, 33.53564, 
    34.03197, 35.69505, 37.58202, 38.97561, 39.48096, 38.97561, 37.58207, 
    35.69675, 34.05672, 33.74171, 55.73597, 57.58053, 59.17378,
  51.26177, 52.61784, 54.62466, 56.08121, 56.40133, 55.91056, 34.71324, 
    35.71807, 37.83025, 40.02993, 41.61595, 42.18832, 41.61595, 40.03, 
    37.8321, 35.74504, 34.94476, 56.85121, 58.95369, 60.79358,
  51.33912, 52.82116, 55.06248, 56.78127, 57.31892, 57.01073, 36.16784, 
    37.62607, 40.05077, 42.44906, 44.1524, 44.76489, 44.1524, 42.44913, 
    40.05275, 37.65419, 36.40941, 58.0087, 60.06858, 61.94059,
  51.36615, 52.90623, 55.27829, 57.18419, 57.92532, 57.83375, 37.2626, 
    39.02143, 41.64272, 44.16174, 45.93305, 46.56796, 45.93305, 44.16182, 
    41.64476, 39.05018, 37.50766, 58.8533, 60.76133, 62.57044,
  51.37195, 52.92738, 55.33902, 57.31044, 58.13225, 58.13365, 37.6586, 
    39.5237, 42.21483, 44.77619, 46.57056, 47.21286, 46.57056, 44.77627, 
    42.2169, 39.55265, 37.90448, 59.15833, 60.99096, 62.76264,
  51.36615, 52.90623, 55.27829, 57.18419, 57.92532, 57.83375, 37.2626, 
    39.02143, 41.64272, 44.16174, 45.93305, 46.56796, 45.93305, 44.16182, 
    41.64476, 39.05018, 37.50766, 58.8533, 60.76133, 62.57044,
  51.33912, 52.82116, 55.06248, 56.78127, 57.31894, 57.0108, 36.16789, 
    37.62613, 40.05084, 42.44913, 44.15248, 44.76497, 44.15248, 42.44921, 
    40.05281, 37.65425, 36.40946, 58.00877, 60.0686, 61.9406,
  51.26177, 52.61785, 54.62469, 56.08138, 56.40192, 55.91195, 34.71474, 
    35.71982, 37.83211, 40.03189, 41.61798, 42.19038, 41.61798, 40.03196, 
    37.83396, 35.74678, 34.94627, 56.85262, 58.9543, 60.7938,
  51.09429, 52.2449, 53.94041, 55.15738, 55.39233, 54.93072, 33.55604, 
    34.05724, 35.72227, 37.6102, 39.00435, 39.5099, 39.00435, 37.61026, 
    35.72398, 34.08199, 33.76215, 55.75041, 57.58681, 59.17617,
  50.81752, 51.70374, 53.07775, 54.18862, 54.58533, 54.44506, 33.46095, 
    33.75732, 34.93229, 36.36831, 37.46109, 37.86045, 37.46109, 36.36837, 
    34.93379, 33.7774, 33.61536, 55.06483, 56.25594, 57.32132,
  50.48119, 51.07206, 52.12305, 53.25059, 54.07667, 54.57817, 54.85091, 
    55.74272, 56.94412, 58.11403, 58.93583, 59.22704, 58.93583, 58.11409, 
    56.94538, 55.75639, 54.94096, 54.95424, 55.14092, 55.41507,
  50.23447, 50.59797, 51.37983, 52.50942, 53.74706, 54.91722, 56.07954, 
    57.5882, 59.03214, 60.14689, 60.81503, 61.03206, 60.81503, 60.14692, 
    59.03278, 57.59488, 56.12304, 55.10995, 54.35389, 53.92636,
  50.10537, 50.32767, 50.91092, 51.98808, 53.49863, 55.22465, 57.12497, 
    59.18222, 60.89444, 62.03902, 62.63302, 62.80716, 62.63302, 62.03904, 
    60.89465, 59.1847, 57.14319, 55.3172, 53.83933, 52.92898,
  50.03724, 50.09667, 50.25145, 50.55619, 51.05235, 51.74329, 52.583, 
    53.40638, 54.0447, 54.45156, 54.65836, 54.71902, 54.65836, 54.4516, 
    54.04498, 53.40813, 52.59147, 51.77579, 51.15349, 50.81635,
  50.10147, 50.2232, 50.50012, 50.96309, 51.60241, 52.37547, 53.25325, 
    54.15094, 54.91011, 55.45541, 55.77, 55.87077, 55.77001, 55.45557, 
    54.91121, 54.15695, 53.27872, 52.46126, 51.83592, 51.48585,
  50.26315, 50.50478, 50.98933, 51.67105, 52.44505, 53.22097, 54.01778, 
    54.92004, 55.78141, 56.48594, 56.94196, 57.09867, 56.94202, 56.4865, 
    55.78502, 54.93802, 54.08716, 53.43301, 52.96425, 52.7058,
  50.57873, 50.97676, 51.67976, 52.50283, 53.25395, 53.85772, 54.38811, 
    55.1591, 56.02582, 56.83331, 57.40824, 57.61634, 57.40842, 56.83486, 
    56.0353, 55.20298, 54.54513, 54.29751, 54.22795, 54.2424,
  51.08964, 51.63134, 52.46805, 53.26596, 53.82541, 54.15916, 54.33606, 
    54.89777, 55.6959, 56.5513, 57.21291, 57.46212, 57.21331, 56.55466, 
    55.71576, 54.98645, 54.63776, 54.94204, 55.39742, 55.78696,
  51.79613, 52.42059, 53.25253, 53.86924, 54.15747, 54.23938, 54.06973, 
    54.3913, 55.07934, 55.96178, 56.70576, 56.99649, 56.70637, 55.96698, 
    55.11138, 54.53948, 54.57603, 55.47485, 56.42672, 57.15817,
  52.65675, 53.33747, 54.10501, 54.47398, 54.43306, 54.19631, 33.24853, 
    33.08464, 33.58711, 34.54715, 35.44409, 35.80567, 35.44464, 34.55243, 
    33.62504, 33.29159, 34.03329, 55.98614, 57.52951, 58.63723,
  53.44526, 54.19617, 54.95351, 55.17693, 54.91646, 54.42946, 33.06484, 
    32.83573, 33.6124, 34.93456, 36.09836, 36.55558, 36.09889, 34.94003, 
    33.65536, 33.0952, 34.11731, 56.73133, 58.80597, 60.23107,
  54.05612, 54.92699, 55.78232, 56.00222, 55.65506, 55.02732, 33.57703, 
    33.62199, 34.77236, 36.38966, 37.73115, 38.24737, 37.73173, 36.39551, 
    34.81861, 33.91068, 34.80477, 57.72489, 60.21687, 61.90279,
  54.45108, 55.45893, 56.47448, 56.79454, 56.48185, 55.85487, 34.57227, 
    34.97535, 36.41684, 38.21957, 39.6634, 40.2126, 39.66403, 38.22584, 
    36.4655, 35.27886, 35.89175, 58.80575, 61.52904, 63.38689,
  54.65524, 55.76894, 56.92804, 57.3675, 57.13507, 56.57741, 35.5008, 
    36.16558, 37.78059, 39.68488, 41.18335, 41.75005, 41.18402, 39.69148, 
    37.83099, 36.47675, 36.85971, 59.65899, 62.4653, 64.41042,
  54.71586, 55.86881, 57.08489, 57.57638, 57.38335, 56.86366, 35.87408, 
    36.63239, 38.30485, 40.24187, 41.75785, 42.33018, 41.75855, 40.2486, 
    38.3559, 36.94601, 37.24345, 59.9843, 62.80538, 64.77554,
  54.65525, 55.76895, 56.92809, 57.36766, 57.13548, 56.57811, 35.50133, 
    36.16612, 37.78116, 39.6855, 41.18401, 41.75074, 41.18469, 39.69211, 
    37.83156, 36.47729, 36.86025, 59.65971, 62.46575, 64.41066,
  54.4511, 55.45905, 56.47493, 56.79596, 56.48519, 55.86071, 34.57745, 
    34.98091, 36.42271, 38.22578, 39.66992, 40.21924, 39.67055, 38.23205, 
    36.47138, 35.28448, 35.89705, 58.81175, 61.53263, 63.38887,
  54.05632, 54.92782, 55.78534, 56.0108, 55.6745, 55.06219, 33.61524, 
    33.66605, 34.81913, 36.43835, 37.78134, 38.29814, 37.78192, 36.44421, 
    34.86546, 33.955, 34.8434, 57.7603, 60.23748, 61.91469,
  53.44653, 54.20076, 54.96851, 55.21639, 55.00167, 54.58267, 33.27469, 
    33.09992, 33.90458, 35.2402, 36.41064, 36.86997, 36.41117, 35.24571, 
    33.94777, 33.36005, 34.3276, 56.88581, 58.896, 60.28601,
  52.66291, 53.35704, 54.16307, 54.61481, 54.71827, 54.69204, 34.0309, 
    34.1336, 34.81722, 35.87402, 36.81203, 37.18423, 36.8126, 35.87937, 
    34.85537, 34.34064, 34.81506, 56.48627, 57.83428, 58.83744,
  51.81974, 52.48702, 53.43084, 54.26391, 54.89277, 55.43259, 55.83005, 
    56.69405, 57.8003, 58.94455, 59.81871, 60.14707, 59.81934, 58.94984, 
    57.83261, 56.84303, 56.34024, 56.68755, 57.23097, 57.73776,
  51.16304, 51.8141, 52.90871, 54.14557, 55.3079, 56.35963, 57.36286, 
    58.79218, 60.32131, 61.68499, 62.6285, 62.96568, 62.62893, 61.68848, 
    60.34185, 58.88426, 57.68071, 57.2057, 57.07237, 57.12805,
  50.76693, 51.39171, 52.57322, 54.09671, 55.65403, 57.06628, 58.45154, 
    60.23279, 62.04999, 63.60077, 64.63518, 64.99678, 64.63538, 63.60254, 
    62.06115, 60.28653, 58.65345, 57.66479, 57.06356, 56.77725,
  50.16629, 50.32495, 50.67499, 51.24941, 52.04582, 53.02829, 54.1585, 
    55.31443, 56.3067, 57.03414, 57.46358, 57.60354, 57.46367, 57.03474, 
    56.3099, 55.32808, 54.20632, 53.16753, 52.38662, 51.95982,
  50.3398, 50.5751, 51.0408, 51.70529, 52.50598, 53.38676, 54.34294, 
    55.35925, 56.28526, 57.02006, 57.4897, 57.65081, 57.49, 57.02187, 
    56.29382, 55.39206, 54.44615, 53.65635, 53.09565, 52.79989,
  50.70573, 51.05361, 51.66663, 52.40619, 53.14262, 53.82332, 54.49094, 
    55.29808, 56.12384, 56.85856, 57.37322, 57.559, 57.37408, 56.86342, 
    56.1452, 55.37406, 54.71145, 54.34981, 54.18375, 54.13791,
  51.29892, 51.73378, 52.41945, 53.11826, 53.6847, 54.11109, 54.45113, 
    55.03385, 55.74071, 56.45146, 56.98937, 57.19099, 56.99141, 56.46228, 
    55.78589, 55.18615, 54.86529, 55.02233, 55.32264, 55.57953,
  52.11533, 52.55264, 53.16952, 53.69522, 54.02983, 54.22044, 54.25826, 
    54.62643, 55.20131, 55.86552, 56.40569, 56.61465, 56.40947, 55.88527, 
    55.28214, 54.89156, 54.94718, 55.62822, 56.33923, 56.84842,
  53.11338, 53.44538, 53.85307, 54.11861, 54.21834, 54.23066, 54.00696, 
    54.16153, 54.58483, 55.19073, 55.73092, 55.94759, 55.73615, 55.21896, 
    54.7048, 54.56584, 55.05038, 56.2254, 57.22841, 57.88319,
  54.26484, 54.43694, 54.57289, 54.5334, 54.3576, 54.13644, 33.28534, 
    32.98101, 33.11538, 33.65234, 34.23136, 34.47625, 34.23615, 33.68159, 
    33.25835, 33.53243, 34.80952, 56.82888, 58.17406, 58.98777,
  55.36643, 55.40287, 55.32443, 55.05319, 54.65739, 54.21807, 32.9653, 
    32.45547, 32.68267, 33.46784, 34.25897, 34.58277, 34.26355, 33.49812, 
    32.84701, 33.15497, 34.99251, 57.58758, 59.28442, 60.25551,
  56.3142, 56.29271, 56.11393, 55.71443, 55.16886, 54.55155, 33.10142, 
    32.68684, 33.17981, 34.21657, 35.16373, 35.53853, 35.16852, 34.2484, 
    33.35735, 33.48055, 35.50702, 58.50171, 60.54819, 61.6893,
  57.01993, 57.01065, 56.83192, 56.40001, 55.78912, 55.08345, 33.66842, 
    33.5034, 34.24526, 35.44523, 36.4758, 36.87552, 36.48093, 35.47869, 
    34.43084, 34.34631, 36.30437, 59.45465, 61.76888, 63.05752,
  57.4436, 57.47506, 57.34063, 56.92612, 56.30478, 55.57975, 34.28289, 
    34.32861, 35.22168, 36.50312, 37.57054, 37.98059, 37.57597, 36.53795, 
    35.41256, 35.19508, 37.03226, 60.19566, 62.66677, 64.05502,
  57.58321, 57.63538, 57.52517, 57.1244, 56.506, 55.78241, 34.54283, 
    34.66644, 35.60824, 36.91356, 37.9911, 38.4039, 37.99665, 36.94893, 
    35.80107, 35.54003, 37.32516, 60.47742, 62.99872, 64.42204,
  57.44367, 57.47531, 57.34139, 56.92804, 56.30864, 55.58563, 34.28751, 
    34.33323, 35.22647, 36.50816, 37.57585, 37.98601, 37.58128, 36.543, 
    35.41738, 35.19982, 37.03712, 60.2019, 62.67115, 64.05795,
  57.02042, 57.01213, 56.8362, 56.41018, 55.80901, 55.11471, 33.69733, 
    33.53432, 34.27735, 35.47852, 36.51021, 36.9104, 36.51535, 35.51202, 
    34.46314, 34.37788, 36.33424, 59.48714, 61.79099, 63.07261,
  56.31678, 56.29972, 56.13263, 55.75653, 55.24895, 54.68042, 33.24557, 
    32.85526, 33.35992, 34.40303, 35.35436, 35.73074, 35.35918, 34.43506, 
    33.53831, 33.65101, 35.6531, 58.63371, 60.63628, 61.75124,
  55.37736, 55.42974, 55.39082, 55.19397, 54.91506, 54.63203, 33.52282, 
    33.16525, 33.4857, 34.31861, 35.13175, 35.46199, 35.13643, 34.34946, 
    33.65186, 33.86725, 35.55023, 58.00955, 59.56919, 60.46468,
  54.30282, 54.5217, 54.76601, 54.91517, 55.01656, 55.15558, 34.80269, 
    34.99603, 35.5206, 36.30356, 37.00593, 37.28685, 37.01088, 36.33334, 
    35.66439, 35.54675, 36.32811, 57.87562, 58.91901, 59.57014,
  53.2233, 53.66764, 54.31596, 54.96009, 55.56062, 56.16656, 56.65408, 
    57.52724, 58.57117, 59.62449, 60.42178, 60.72068, 60.4272, 59.6534, 
    58.69301, 57.93768, 57.72285, 58.24975, 58.8026, 59.21315,
  52.38347, 53.04214, 54.0922, 55.21878, 56.24533, 57.16156, 57.99543, 
    59.25325, 60.66041, 61.98075, 62.93198, 63.27985, 62.93606, 62.00184, 
    60.74667, 59.53949, 58.75851, 58.78556, 59.06317, 59.34851,
  51.85759, 52.65284, 53.97689, 55.43748, 56.73684, 57.81356, 58.80541, 
    60.24273, 61.8437, 63.33821, 64.41232, 64.80454, 64.41477, 63.3515, 
    61.90091, 60.4438, 59.38137, 59.15823, 59.30833, 59.53761,
  50.51148, 50.80848, 51.39492, 52.23613, 53.26495, 54.41767, 55.68222, 
    57.01475, 58.23996, 59.224, 59.85963, 60.07918, 59.86066, 59.22888, 
    58.25892, 57.07674, 55.85416, 54.82568, 54.09838, 53.71603,
  50.83932, 51.17644, 51.79211, 52.59027, 53.47702, 54.40306, 55.38178, 
    56.45279, 57.47076, 58.32044, 58.88903, 59.08985, 58.8915, 58.33123, 
    57.50901, 56.56708, 55.67094, 55.02715, 54.63358, 54.45531,
  51.45231, 51.81763, 52.42332, 53.10704, 53.76164, 54.36647, 54.95014, 
    55.68181, 56.43952, 57.12503, 57.61324, 57.79202, 57.61887, 57.1483, 
    56.51725, 55.89928, 55.45989, 55.37258, 55.44788, 55.55311,
  52.31684, 52.63807, 53.12658, 53.60941, 54.00349, 54.31679, 54.54414, 
    54.98609, 55.52175, 56.06588, 56.48283, 56.64184, 56.49384, 56.10979, 
    55.66273, 55.36242, 55.37357, 55.82763, 56.3123, 56.65158,
  53.36435, 53.54244, 53.79432, 54.01417, 54.16604, 54.26677, 54.21976, 
    54.4352, 54.78613, 55.20855, 55.56225, 55.70366, 55.58028, 55.27971, 
    55.01139, 55.02156, 55.45476, 56.35978, 57.10608, 57.56968,
  54.52518, 54.47295, 54.39748, 54.32365, 54.26527, 54.22314, 53.96201, 
    53.97697, 54.1448, 54.44445, 54.7365, 54.86118, 54.76009, 54.54082, 
    54.45993, 54.81071, 55.68488, 56.95015, 57.81515, 58.29831,
  55.80982, 55.48405, 55.03281, 54.62724, 54.3199, 54.08689, 33.30638, 
    32.9014, 32.7192, 32.82909, 33.05349, 33.16479, 33.07587, 32.93135, 
    33.09759, 34.01219, 35.68684, 57.55593, 58.56593, 59.08259,
  57.07093, 56.49318, 55.70597, 55.00968, 54.47454, 54.0402, 32.89268, 
    32.19736, 31.94157, 32.16484, 32.53138, 32.70099, 32.5528, 32.27251, 
    32.3855, 33.61453, 36.00393, 58.25109, 59.43945, 60.0079,
  58.23342, 57.46326, 56.42039, 55.49509, 54.76036, 54.12223, 32.7074, 
    31.94285, 31.81361, 32.22411, 32.72484, 32.94044, 32.74669, 32.33651, 
    32.29928, 33.58224, 36.42748, 59.01534, 60.43153, 61.08603,
  59.17924, 58.28643, 57.08063, 56.00394, 55.12811, 54.33922, 32.83677, 
    32.19231, 32.25064, 32.80635, 33.38412, 33.62265, 33.40685, 32.92248, 
    32.75806, 33.95845, 36.97525, 59.76834, 61.39527, 62.13982,
  59.79781, 58.84376, 57.55594, 56.39936, 55.44569, 54.5752, 33.09019, 
    32.59185, 32.7821, 33.41299, 34.0224, 34.26908, 34.04599, 33.53214, 
    33.30111, 34.41864, 37.45905, 60.33877, 62.10853, 62.91953,
  60.01308, 59.04175, 57.73074, 56.551, 55.57458, 54.68092, 33.21476, 
    32.77591, 33.01062, 33.66328, 34.28055, 34.52901, 34.3045, 33.78367, 
    33.5336, 34.62065, 37.65575, 60.55756, 62.37625, 63.2107,
  59.79873, 58.84591, 57.5611, 56.41001, 55.46418, 54.60142, 33.11196, 
    32.61355, 32.80403, 33.43546, 34.04551, 34.29247, 34.06911, 33.55473, 
    33.32348, 34.44144, 37.4823, 60.36697, 62.13027, 62.93629,
  59.18354, 58.29578, 57.10183, 56.04606, 55.20027, 54.44452, 32.9385, 
    32.30233, 32.36444, 32.92243, 33.5022, 33.74159, 33.52503, 33.03909, 
    32.8737, 34.07231, 37.08083, 59.87924, 61.47871, 62.20506,
  58.24984, 57.49626, 56.49079, 55.6291, 54.98521, 54.45634, 33.08912, 
    32.39678, 32.30714, 32.73599, 33.24563, 33.46418, 33.26789, 32.85016, 
    32.79778, 34.04335, 36.81365, 59.3628, 60.69072, 61.29353,
  57.1238, 56.5915, 55.9023, 55.36452, 55.04884, 54.88615, 34.01264, 
    33.62982, 33.59814, 33.95049, 34.37878, 34.56649, 34.40117, 34.06145, 
    34.04826, 35.04977, 37.12389, 59.13324, 60.11214, 60.56691,
  55.95485, 55.73318, 55.49392, 55.40709, 55.51154, 55.76835, 35.67435, 
    35.98938, 36.43411, 36.99328, 37.4731, 37.66562, 37.49636, 37.09752, 
    36.81382, 37.09931, 38.0793, 59.34394, 60.01166, 60.34951,
  54.86639, 55.01185, 55.31141, 55.74866, 56.28367, 56.88136, 57.37397, 
    58.18143, 59.08951, 59.9754, 60.6355, 60.88482, 60.6603, 60.07526, 
    59.41396, 59.04525, 59.19634, 59.87193, 60.38696, 60.69653,
  54.05888, 54.5465, 55.33808, 56.20927, 57.02217, 57.75657, 58.38668, 
    59.39997, 60.55285, 61.65902, 62.4707, 62.77325, 62.49074, 61.73768, 
    60.80347, 60.06704, 59.84655, 60.37186, 60.96632, 61.39151,
  53.55615, 54.27588, 55.39585, 56.53548, 57.48664, 58.25213, 58.91021, 
    59.9889, 61.24635, 62.46982, 63.37572, 63.71347, 63.38984, 62.52729, 
    61.43724, 60.52259, 60.15197, 60.65055, 61.36932, 61.92135,
  51.71099, 52.16344, 52.97528, 54.00272, 55.11381, 56.24301, 57.4129, 
    58.68287, 59.90969, 60.95821, 61.67509, 61.93341, 61.6881, 61.0028, 
    60.03556, 58.9921, 58.07666, 57.49457, 57.1951, 57.08311,
  52.21804, 52.58825, 53.24149, 54.05559, 54.93139, 55.82517, 56.74224, 
    57.77122, 58.76793, 59.61837, 60.19922, 60.41081, 60.22153, 59.6904, 
    58.95785, 58.20549, 57.6061, 57.33024, 57.24728, 57.25138,
  53.06678, 53.28548, 53.67151, 54.15617, 54.68622, 55.23613, 55.76817, 
    56.43524, 57.09278, 57.6609, 58.05432, 58.20384, 58.09367, 57.78287, 
    57.39812, 57.09093, 56.97661, 57.16164, 57.37735, 57.53245,
  54.11395, 54.12758, 54.1861, 54.31358, 54.50505, 54.73561, 54.89395, 
    55.21172, 55.54275, 55.84564, 56.06836, 56.16447, 56.13208, 56.0386, 
    56.00975, 56.16894, 56.55081, 57.17299, 57.6227, 57.88021,
  55.23177, 55.01565, 54.73017, 54.51948, 54.42819, 54.41969, 54.2877, 
    54.32802, 54.3929, 54.48163, 54.56976, 54.62642, 54.66169, 54.75854, 
    55.0537, 55.64392, 56.45757, 57.39861, 57.95793, 58.24225,
  56.35295, 55.90314, 55.27515, 54.74697, 54.41914, 54.24029, 53.89733, 
    53.71453, 53.54533, 53.43851, 53.40211, 53.42096, 53.51694, 53.79401, 
    54.41113, 55.43568, 56.64194, 57.76726, 58.32276, 58.56846,
  57.5442, 56.85347, 55.86098, 54.98139, 54.38153, 54.00209, 33.22703, 
    32.66119, 32.0947, 31.67269, 31.44457, 31.39896, 31.55993, 32.06456, 
    33.14132, 34.86591, 36.7344, 58.17286, 58.72622, 58.94181,
  58.72708, 57.80729, 56.46352, 55.24102, 54.36764, 53.76731, 32.66022, 
    31.74258, 30.92183, 30.41754, 30.20989, 30.18349, 30.32441, 30.84676, 
    32.18187, 34.53379, 37.07624, 58.59418, 59.16938, 59.36737,
  59.86562, 58.73379, 57.06229, 55.51486, 54.36945, 53.52375, 32.08621, 
    30.91912, 30.01719, 29.57664, 29.46108, 29.47278, 29.57626, 30.03029, 
    31.43513, 34.20753, 37.33709, 58.99234, 59.6408, 59.84745,
  60.84163, 59.53119, 57.58617, 55.77038, 54.39863, 53.33825, 31.66487, 
    30.42572, 29.59266, 29.27104, 29.24243, 29.28381, 29.35819, 29.73489, 
    31.0957, 34.05011, 37.56765, 59.34817, 60.08515, 60.31063,
  61.51002, 60.07864, 57.95137, 55.96088, 54.44427, 53.2446, 31.44696, 
    30.23807, 29.50079, 29.26582, 29.28592, 29.34219, 29.40258, 29.73413, 
    31.04122, 34.04203, 37.75515, 59.61404, 60.41758, 60.65795,
  61.75113, 60.27847, 58.09074, 56.04537, 54.48629, 53.24528, 31.40689, 
    30.2217, 29.52337, 29.31732, 29.35186, 29.41236, 29.46912, 29.78758, 
    31.07545, 34.08271, 37.85326, 59.7432, 60.5669, 60.8094,
  61.52253, 60.09923, 57.98873, 56.02373, 54.53891, 53.36994, 31.56073, 
    30.35436, 29.61712, 29.38122, 29.401, 29.4574, 29.51832, 29.85192, 
    31.16348, 34.16732, 37.87694, 59.75179, 60.53497, 60.76078,
  60.88361, 59.59718, 57.70121, 55.95921, 54.68065, 53.71948, 32.05722, 
    30.86393, 30.05369, 29.73825, 29.71069, 29.75269, 29.82881, 30.20975, 
    31.57248, 34.50639, 37.97388, 59.76175, 60.43435, 60.61972,
  59.98167, 58.90656, 57.3485, 55.96783, 55.03248, 54.42551, 33.14168, 
    32.20166, 31.45828, 31.10066, 31.01999, 31.04212, 31.14072, 31.56918, 
    32.89772, 35.50241, 38.40642, 59.97201, 60.47363, 60.5991,
  59.00753, 58.2007, 57.07584, 56.16227, 55.66548, 55.49561, 34.87653, 
    34.55103, 34.23838, 34.08781, 34.07543, 34.11172, 34.19734, 34.53143, 
    35.5073, 37.3362, 39.33324, 60.51489, 60.85544, 60.93526,
  58.14005, 57.6367, 56.99146, 56.57162, 56.49524, 56.68351, 36.7188, 
    37.04644, 37.3408, 37.62168, 37.84649, 37.95732, 37.96623, 38.02007, 
    38.39471, 39.29259, 40.42277, 61.28375, 61.61273, 61.73042,
  57.46865, 57.27084, 57.0848, 57.09578, 57.32619, 57.69824, 58.00933, 
    58.54484, 59.09657, 59.60995, 59.99293, 60.16171, 60.11611, 59.98861, 
    60.02422, 60.43527, 61.16311, 62.01968, 62.53558, 62.79817,
  57.08607, 57.13111, 57.27657, 57.54579, 57.89996, 58.28689, 58.57641, 
    59.15222, 59.79057, 60.40102, 60.85803, 61.05129, 60.96547, 60.7272, 
    60.58741, 60.80399, 61.45341, 62.51916, 63.33596, 63.81101,
  56.8821, 57.07542, 57.40727, 57.80011, 58.19167, 58.55635, 58.81178, 
    59.3804, 60.03593, 60.67422, 61.15439, 61.35206, 61.24266, 60.94907, 
    60.73021, 60.87807, 61.5402, 62.76635, 63.80371, 64.42829,
  53.06672, 53.50178, 54.26387, 55.19836, 56.17712, 57.14322, 58.11366, 
    59.18063, 60.21093, 61.0934, 61.70066, 61.92776, 61.74492, 61.22438, 
    60.52735, 59.85254, 59.37413, 59.24421, 59.3037, 59.39441,
  53.56145, 53.85746, 54.39423, 55.08619, 55.85137, 56.64074, 57.43369, 
    58.33318, 59.19576, 59.92682, 60.42772, 60.62136, 60.49275, 60.11037, 
    59.61428, 59.1678, 58.89887, 58.92444, 59.04293, 59.14671,
  54.36001, 54.44196, 54.63431, 54.95434, 55.38306, 55.87968, 56.36032, 
    56.96545, 57.54016, 58.02084, 58.35139, 58.49306, 58.45193, 58.29449, 
    58.1334, 58.07623, 58.16893, 58.46902, 58.69852, 58.83578,
  55.30853, 55.1613, 54.9873, 54.91315, 54.98211, 55.15813, 55.28085, 
    55.54312, 55.78451, 55.98292, 56.12707, 56.21515, 56.27534, 56.37767, 
    56.61062, 57.01511, 57.52715, 58.12809, 58.46822, 58.63742,
  56.28649, 55.93502, 55.43058, 54.99894, 54.7445, 54.63834, 54.44473, 
    54.39334, 54.32595, 54.26596, 54.24308, 54.28621, 54.4445, 54.79887, 
    55.42163, 56.28122, 57.18129, 58.01591, 58.41469, 58.58975,
  57.23615, 56.71328, 55.92139, 55.17257, 54.6382, 54.3047, 53.86946, 
    53.55463, 53.21204, 52.91376, 52.73358, 52.73174, 52.98042, 53.58022, 
    54.59613, 55.90775, 57.14443, 58.09024, 58.47351, 58.61588,
  58.22968, 57.54188, 56.45768, 55.36963, 54.5301, 53.95428, 33.1013, 
    32.39922, 31.63955, 30.97462, 30.54616, 30.45638, 30.80429, 31.72628, 
    33.30999, 35.32424, 37.0837, 58.23539, 58.59274, 58.70354,
  59.20323, 58.36004, 56.99419, 55.5729, 54.42655, 53.59201, 32.39954, 
    31.31819, 30.22876, 29.37332, 28.88071, 28.77974, 29.14662, 30.22028, 
    32.2579, 34.96801, 37.27113, 58.38203, 58.72348, 58.80658,
  60.132, 59.13862, 57.49965, 55.75294, 54.29885, 53.1842, 31.6293, 30.2217, 
    28.9395, 28.05538, 27.61075, 27.53645, 27.88084, 28.96822, 31.26292, 
    34.53192, 37.35231, 58.48847, 58.84936, 58.92085,
  60.92307, 59.79798, 57.92246, 55.89788, 54.181, 52.81659, 30.95424, 
    29.36505, 28.06084, 27.26167, 26.90632, 26.8656, 27.17541, 28.20169, 
    30.56451, 34.169, 37.38179, 58.57167, 58.96827, 59.03636,
  61.4645, 60.24888, 58.21324, 56.00468, 54.11655, 52.5859, 30.52327, 
    28.88029, 27.63097, 26.92215, 26.6319, 26.61278, 26.89955, 27.86975, 
    30.21995, 33.97383, 37.41626, 58.65261, 59.07813, 59.14408,
  61.66739, 60.42373, 58.33989, 56.07922, 54.14627, 52.5709, 30.43325, 
    28.785, 27.56467, 26.889, 26.61972, 26.60738, 26.88765, 27.84025, 
    30.18223, 33.97769, 37.49325, 58.75691, 59.18633, 59.24628,
  61.50809, 60.31048, 58.3102, 56.15205, 54.32389, 52.85236, 30.77985, 
    29.15063, 27.90464, 27.19204, 26.89798, 26.87823, 27.16917, 28.14992, 
    30.51221, 34.26448, 37.68927, 58.95135, 59.34592, 59.39132,
  61.0496, 59.97057, 58.18478, 56.28748, 54.72403, 53.52314, 31.70923, 
    30.22859, 28.98979, 28.21315, 27.86093, 27.82198, 28.14007, 29.17833, 
    31.52886, 35.06039, 38.16439, 59.36286, 59.67688, 59.69675,
  60.43183, 59.52936, 58.06488, 56.56152, 55.3998, 54.61152, 33.31329, 
    32.281, 31.29918, 30.59966, 30.24328, 30.19807, 30.5303, 31.54505, 
    33.64847, 36.59706, 39.084, 60.11298, 60.3244, 60.31917,
  59.83056, 59.13606, 58.04876, 57.00311, 56.29408, 55.9441, 35.33863, 
    34.98521, 34.57324, 34.24076, 34.06525, 34.07334, 34.3469, 35.10776, 
    36.60305, 38.6453, 40.36872, 61.16427, 61.33429, 61.34235,
  59.39717, 58.9055, 58.17713, 57.54591, 57.20814, 57.15946, 37.07437, 
    37.24743, 37.36745, 37.46255, 37.55217, 37.64879, 37.81915, 38.22953, 
    39.07691, 40.33133, 41.52711, 62.25424, 62.5449, 62.65096,
  59.17273, 58.84331, 58.39238, 58.05968, 57.95165, 58.03087, 58.10472, 
    58.36728, 58.62297, 58.85822, 59.05209, 59.19049, 59.32203, 59.58945, 
    60.17145, 61.10884, 62.16418, 63.11312, 63.66266, 63.93203,
  59.17069, 58.92442, 58.60876, 58.4057, 58.37215, 58.45867, 58.48354, 
    58.74444, 59.02555, 59.29556, 59.51658, 59.65973, 59.76157, 59.95632, 
    60.4333, 61.29375, 62.40836, 63.65327, 64.47883, 64.91586,
  59.21523, 58.99483, 58.72338, 58.56289, 58.55022, 58.62914, 58.62217, 
    58.86477, 59.13332, 59.39254, 59.60334, 59.73462, 59.81862, 59.9856, 
    60.43401, 61.29945, 62.49789, 63.92664, 64.91972, 65.45065,
  55.81309, 56.01311, 56.38552, 56.87995, 57.4357, 58.00378, 58.5521, 
    59.17956, 59.75864, 60.23639, 60.56966, 60.73323, 60.74551, 60.68098, 
    60.65385, 60.76787, 61.06504, 61.58159, 62.05217, 62.33811,
  56.05602, 56.14833, 56.3535, 56.68021, 57.1029, 57.57658, 58.03752, 
    58.59618, 59.11361, 59.54184, 59.84714, 60.01388, 60.06663, 60.07791, 
    60.14489, 60.33697, 60.65805, 61.1385, 61.51971, 61.74054,
  56.45506, 56.38807, 56.33363, 56.38, 56.55856, 56.83999, 57.11081, 
    57.51004, 57.88176, 58.19128, 58.4249, 58.58698, 58.71422, 58.87451, 
    59.13285, 59.49863, 59.91114, 60.39041, 60.67673, 60.8241,
  56.9578, 56.73405, 56.40499, 56.12349, 55.98308, 55.98515, 55.97068, 
    56.10976, 56.23795, 56.34687, 56.45544, 56.59948, 56.83409, 57.21919, 
    57.77206, 58.41946, 59.0152, 59.55861, 59.79861, 59.90146,
  57.50723, 57.16044, 56.59442, 55.99689, 55.51732, 55.19997, 54.86443, 
    54.68257, 54.50224, 54.35266, 54.29626, 54.41013, 54.77423, 55.43982, 
    56.36377, 57.36849, 58.20502, 58.83844, 59.07341, 59.15837,
  58.04918, 57.61788, 56.86795, 55.99575, 55.19884, 54.57247, 53.94614, 
    53.43553, 52.92987, 52.49879, 52.25561, 52.32759, 52.82962, 53.81214, 
    55.16057, 56.55759, 57.63089, 58.29862, 58.52578, 58.59373,
  58.62006, 58.11685, 57.1962, 56.05162, 54.93196, 53.99482, 32.93413, 
    31.98766, 31.03864, 30.2012, 29.66418, 29.63739, 30.29928, 31.72065, 
    33.69505, 35.67754, 37.08512, 57.8992, 58.11396, 58.16682,
  59.14889, 58.58871, 57.52241, 56.13029, 54.70101, 53.44712, 31.9866, 
    30.59444, 29.23133, 28.07337, 27.34995, 27.27148, 28.04872, 29.85092, 
    32.45931, 35.05985, 36.82324, 57.55682, 57.76265, 57.80143,
  59.62109, 59.01148, 57.81445, 56.19231, 54.46432, 52.89012, 31.02143, 
    29.21542, 27.53374, 26.20548, 25.4334, 25.35285, 26.17066, 28.18941, 
    31.28796, 34.44212, 36.55253, 57.23932, 57.44979, 57.48077,
  60.00298, 59.35442, 58.05219, 56.24087, 54.26105, 52.4065, 30.16241, 
    28.0395, 26.19309, 24.85508, 24.13881, 24.08465, 24.88395, 26.9552, 
    30.33845, 33.90688, 36.30716, 56.99175, 57.21376, 57.23972,
  60.26802, 59.59804, 58.23387, 56.30628, 54.1672, 52.1285, 29.60889, 
    27.30637, 25.41923, 24.13962, 23.49455, 23.46564, 24.23544, 26.28734, 
    29.79095, 33.60128, 36.19197, 56.89927, 57.12983, 57.15068,
  60.40734, 59.74085, 58.37561, 56.43505, 54.27176, 52.1993, 29.57611, 
    27.22813, 25.34222, 24.08888, 23.46803, 23.44819, 24.21195, 26.26065, 
    29.80145, 33.68507, 36.3313, 57.06798, 57.29219, 57.30506,
  60.44458, 59.81179, 58.51757, 56.68534, 54.65809, 52.73804, 30.24677, 
    28.01793, 26.16948, 24.89425, 24.24149, 24.21416, 25.00475, 27.0857, 
    30.58682, 34.34533, 36.87043, 57.61794, 57.81243, 57.8135,
  60.44323, 59.87354, 58.71913, 57.1091, 55.36757, 53.77694, 31.69482, 
    29.84813, 28.21367, 26.99276, 26.3236, 26.29242, 27.11053, 29.15754, 
    32.40204, 35.74308, 37.935, 58.63996, 58.78988, 58.78187,
  60.4945, 60.00442, 59.0299, 57.7085, 56.33586, 55.16307, 33.70132, 
    32.48169, 31.34126, 30.42238, 29.89245, 29.90332, 30.6681, 32.44128, 
    35.08926, 37.74012, 39.46946, 60.08383, 60.21782, 60.22316,
  60.68135, 60.25908, 59.44795, 58.39739, 57.36585, 56.55524, 35.70121, 
    35.08308, 34.50084, 34.01836, 33.75505, 33.84833, 34.47536, 35.80949, 
    37.75274, 39.73915, 41.1156, 61.68386, 61.89042, 61.95463,
  61.03311, 60.6333, 59.90754, 59.02813, 58.21645, 57.61449, 37.09736, 
    36.83003, 36.599, 36.41983, 36.36193, 36.51907, 37.02363, 38.01482, 
    39.47697, 41.09114, 42.38546, 63.08098, 63.46316, 63.63334,
  61.47578, 61.04222, 60.30937, 59.49283, 58.78551, 58.26579, 57.8411, 
    57.60825, 57.41539, 57.28328, 57.26842, 57.44691, 57.92765, 58.82578, 
    60.14809, 61.67973, 63.05485, 64.06815, 64.66346, 64.94741,
  61.93606, 61.41727, 60.59007, 59.73626, 59.04425, 58.54624, 58.08197, 
    57.85164, 57.65711, 57.52074, 57.5002, 57.66822, 58.12796, 58.99592, 
    60.30547, 61.88694, 63.39494, 64.68275, 65.43501, 65.79809,
  62.24185, 61.64143, 60.71829, 59.81538, 59.12431, 58.64305, 58.1643, 
    57.92628, 57.71051, 57.54432, 57.49446, 57.63959, 58.08596, 58.95707, 
    60.30274, 61.96421, 63.58045, 65.00711, 65.82761, 66.21728,
  57.86327, 57.84065, 57.84573, 57.92899, 58.0965, 58.31416, 58.51968, 
    58.81176, 59.06806, 59.27435, 59.44236, 59.59886, 59.79338, 60.09554, 
    60.56742, 61.2149, 61.96605, 62.79242, 63.41161, 63.75004,
  57.86126, 57.80251, 57.74225, 57.74558, 57.83673, 57.99487, 58.14604, 
    58.40931, 58.65276, 58.85983, 59.04008, 59.21915, 59.445, 59.78073, 
    60.27185, 60.90214, 61.58858, 62.32305, 62.83867, 63.11591,
  57.88388, 57.76017, 57.57882, 57.42744, 57.36278, 57.39047, 57.41499, 
    57.59043, 57.7704, 57.94002, 58.11183, 58.31587, 58.60058, 59.01667, 
    59.57766, 60.22666, 60.85635, 61.48326, 61.85791, 62.04948,
  57.97282, 57.77304, 57.43942, 57.07508, 56.77424, 56.58218, 56.39033, 
    56.38116, 56.40524, 56.46033, 56.57394, 56.79212, 57.16889, 57.73566, 
    58.45598, 59.21262, 59.85806, 60.41878, 60.68086, 60.80087,
  58.13091, 57.86259, 57.37817, 56.77958, 56.19239, 55.70882, 55.23663, 
    54.9444, 54.71078, 54.56015, 54.55187, 54.76513, 55.26875, 56.06855, 
    57.05585, 58.02716, 58.77801, 59.3187, 59.52483, 59.60455,
  58.31559, 57.99983, 57.3942, 56.58091, 55.70447, 54.90434, 54.14208, 
    53.50327, 52.9431, 52.5186, 52.33493, 52.52361, 53.18421, 54.29585, 
    55.64789, 56.91068, 57.81325, 58.32706, 58.51362, 58.57374,
  58.54284, 58.18931, 57.47539, 56.45467, 55.28756, 54.16419, 32.96343, 
    31.84648, 30.83185, 30.00129, 29.52567, 29.63249, 30.49521, 32.0761, 
    34.00227, 35.72404, 36.86339, 57.50769, 57.69267, 57.74588,
  58.73915, 58.36648, 57.57742, 56.38559, 54.95041, 53.50047, 31.84537, 
    30.21168, 28.72217, 27.49782, 26.76645, 26.81311, 27.88297, 29.97319, 
    32.54959, 34.78754, 36.20697, 56.8195, 57.01894, 57.07378,
  58.89881, 58.51877, 57.67734, 56.34285, 54.66341, 52.8988, 30.81104, 
    28.70041, 26.81795, 25.32943, 24.46991, 24.4968, 25.6904, 28.15231, 
    31.28328, 33.99427, 35.67833, 56.25601, 56.47638, 56.53735,
  59.02387, 58.64562, 57.77457, 56.33624, 54.46201, 52.4325, 29.9543, 
    27.44941, 25.3058, 23.71626, 22.85674, 22.89685, 24.12317, 26.77534, 
    30.29561, 33.38531, 35.28974, 55.8672, 56.10695, 56.17307,
  59.13706, 58.76879, 57.89394, 56.40578, 54.41962, 52.22537, 29.45771, 
    26.69984, 24.43369, 22.84673, 22.03639, 22.09713, 23.31474, 26.03178, 
    29.76583, 33.09612, 35.14691, 55.75344, 56.0049, 56.07262,
  59.27582, 58.92602, 58.07758, 56.60905, 54.62678, 52.42107, 29.55882, 
    26.74596, 24.46298, 22.88933, 22.09861, 22.16988, 23.3928, 26.13596, 
    29.93252, 33.32343, 35.40266, 56.0452, 56.29245, 56.35664,
  59.49195, 59.16867, 58.37753, 57.00313, 55.15383, 53.11669, 30.43758, 
    27.83808, 25.6787, 24.13649, 23.33615, 23.41152, 24.66107, 27.38585, 
    31.05086, 34.26236, 36.20861, 56.86075, 57.08581, 57.14357,
  59.84539, 59.55112, 58.83624, 57.61071, 55.99461, 54.26833, 32.05279, 
    29.96569, 28.18033, 26.83527, 26.10733, 26.20894, 27.43335, 29.94931, 
    33.1767, 35.94212, 37.60811, 58.22012, 58.42387, 58.48258,
  60.38121, 60.10332, 59.45248, 58.37959, 57.02029, 55.63675, 34.01442, 
    32.57048, 31.3423, 30.40055, 29.9023, 30.06966, 31.15127, 33.21936, 
    35.78987, 38.00888, 39.39093, 59.94901, 60.17354, 60.257,
  61.09401, 60.79852, 60.15801, 59.17876, 58.01234, 56.88711, 35.7577, 
    34.8195, 34.06285, 33.50827, 33.26181, 33.49447, 34.39278, 36.00717, 
    38.02377, 39.86721, 41.1356, 61.70702, 62.02233, 62.16208,
  61.90918, 61.54914, 60.84014, 59.85872, 58.77562, 57.78011, 36.8903, 
    36.23861, 35.7455, 35.41157, 35.31419, 35.57938, 36.34835, 37.68013, 
    39.40036, 41.11699, 42.45861, 63.1686, 63.62757, 63.84517,
  62.68224, 62.22569, 61.39454, 60.34499, 59.26847, 58.31283, 57.5008, 
    56.90801, 56.44357, 56.13546, 56.06511, 56.34471, 57.09196, 58.35671, 
    60.01085, 61.73825, 63.19016, 64.18448, 64.79447, 65.08667,
  63.32349, 62.75589, 61.77201, 60.61099, 59.49648, 58.54961, 57.70433, 
    57.14006, 56.68604, 56.37634, 56.29963, 56.56887, 57.30191, 58.56019, 
    60.24337, 62.0512, 63.61521, 64.83569, 65.53839, 65.87393,
  63.71025, 63.06009, 61.96071, 60.71386, 59.57031, 58.63237, 57.77563, 
    57.21798, 56.75327, 56.41984, 56.31654, 56.56498, 57.29214, 58.5733, 
    60.31945, 62.21717, 63.86414, 65.18712, 65.92061, 66.26506,
  59.82101, 59.60434, 59.26799, 58.9338, 58.67252, 58.4871, 58.31425, 
    58.26622, 58.2294, 58.21775, 58.28085, 58.48117, 58.88572, 59.54612, 
    60.45987, 61.53405, 62.60637, 63.62276, 64.31503, 64.6731,
  59.60248, 59.41198, 59.10285, 58.77233, 58.48906, 58.27328, 58.0677, 
    58.01262, 57.98898, 58.0052, 58.10217, 58.33379, 58.7577, 59.4131, 
    60.28423, 61.27557, 62.24117, 63.1591, 63.76925, 64.08636,
  59.27347, 59.10378, 58.80723, 58.45266, 58.10906, 57.82301, 57.54063, 
    57.44419, 57.4085, 57.43828, 57.56628, 57.83806, 58.29912, 58.96784, 
    59.80333, 60.69947, 61.52521, 62.2984, 62.77494, 63.02118,
  58.94046, 58.77093, 58.44939, 58.01952, 57.55342, 57.12906, 56.70504, 
    56.49171, 56.37447, 56.36262, 56.48843, 56.79626, 57.32073, 58.05133, 
    58.90754, 59.75916, 60.4783, 61.10467, 61.44166, 61.61,
  58.66475, 58.47744, 58.09803, 57.54649, 56.89659, 56.25743, 55.62836, 
    55.19321, 54.88983, 54.74557, 54.80807, 55.13681, 55.76272, 56.63673, 
    57.61585, 58.52225, 59.21548, 59.72043, 59.95554, 60.0633,
  58.44038, 58.23442, 57.79369, 57.10893, 56.24689, 55.34165, 54.46988, 
    53.70699, 53.1109, 52.73719, 52.66646, 52.9982, 53.77533, 54.8975, 
    56.11996, 57.18235, 57.92733, 58.32943, 58.51526, 58.58988,
  58.29145, 58.06732, 57.56483, 56.74267, 55.65755, 54.4649, 33.18476, 
    31.91899, 30.87245, 30.12051, 29.79332, 30.08251, 31.08945, 32.64782, 
    34.32632, 35.70519, 36.60004, 57.10398, 57.28426, 57.35058,
  58.15764, 57.93209, 57.39786, 56.472, 55.18406, 53.69356, 31.92031, 
    30.06279, 28.47464, 27.2692, 26.64346, 26.89311, 28.19932, 30.32729, 
    32.59764, 34.3914, 35.524, 56.07909, 56.29483, 56.37453,
  58.04347, 57.82951, 57.28839, 56.29129, 54.83229, 53.06784, 30.85222, 
    28.44921, 26.38557, 24.82086, 23.98688, 24.21553, 25.7549, 28.37447, 
    31.19294, 33.37986, 34.73693, 55.30376, 55.5626, 55.66249,
  57.97372, 57.78022, 57.2532, 56.22116, 54.64162, 52.6626, 30.0722, 
    27.21151, 24.78831, 23.01457, 22.10171, 22.33472, 24.00202, 26.95574, 
    30.2031, 32.71119, 34.24579, 54.83673, 55.13041, 55.24732,
  58.0015, 57.83257, 57.33513, 56.30608, 54.67429, 52.57851, 29.72426, 
    26.56377, 23.93363, 22.08248, 21.17205, 21.42116, 23.13915, 26.26949, 
    29.78123, 32.49492, 34.13878, 54.77532, 55.09006, 55.2175,
  58.19333, 58.04839, 57.58998, 56.60128, 54.9998, 52.92238, 30.01196, 
    26.81565, 24.16668, 22.32061, 21.42596, 21.69175, 23.4356, 26.61506, 
    30.18035, 32.91848, 34.56308, 55.24022, 55.55772, 55.68869,
  58.61531, 58.48721, 58.06625, 57.14386, 55.64848, 53.72758, 31.04102, 
    28.15132, 25.73986, 24.02465, 23.18267, 23.47379, 25.2025, 28.24836, 
    31.58135, 34.11081, 35.62574, 56.30241, 56.60883, 56.74049,
  59.31101, 59.18146, 58.77529, 57.91467, 56.55868, 54.87172, 32.63572, 
    30.31866, 28.40401, 27.03122, 26.37348, 26.71349, 28.30381, 30.95211, 
    33.77748, 35.93181, 37.25154, 57.88223, 58.18639, 58.32568,
  60.26823, 60.10477, 59.66351, 58.81786, 57.56985, 56.09492, 34.34842, 
    32.61843, 31.2512, 30.31175, 29.92409, 30.31838, 31.67369, 33.81295, 
    36.09941, 37.92525, 39.12506, 59.71581, 60.05482, 60.21801,
  61.39417, 61.15689, 60.61493, 59.70963, 58.49246, 57.14145, 35.74747, 
    34.43192, 33.45292, 32.83108, 32.64817, 33.06858, 34.2183, 35.98227, 
    37.9361, 39.62961, 40.85883, 61.46893, 61.88369, 62.0864,
  62.53421, 62.19237, 61.49549, 60.46119, 59.19428, 57.876, 36.63226, 
    35.57378, 34.81686, 34.3642, 34.28506, 34.70677, 35.73089, 37.29906, 
    39.12517, 40.84122, 42.18908, 62.89484, 63.40485, 63.65515,
  63.51184, 63.06408, 62.2049, 61.02201, 59.66784, 58.3252, 57.13622, 
    56.18536, 55.48036, 55.05846, 55.00574, 55.43839, 56.44009, 57.96301, 
    59.77145, 61.53004, 62.95934, 63.8902, 64.50016, 64.79883,
  64.24919, 63.7085, 62.70017, 61.37117, 59.92336, 58.55061, 57.31762, 
    56.42261, 55.75093, 55.34234, 55.29246, 55.72145, 56.71927, 58.25515, 
    60.11107, 61.94259, 63.44072, 64.55519, 65.22014, 65.54564,
  64.66946, 64.07263, 62.96925, 61.54223, 60.03004, 58.63708, 57.38112, 
    56.50455, 55.8376, 55.41885, 55.35266, 55.77018, 56.77525, 58.35064, 
    60.27633, 62.18048, 63.72656, 64.92026, 65.60181, 65.93331,
  62.2062, 61.8273, 61.15392, 60.31736, 59.4449, 58.62641, 57.86473, 
    57.33231, 56.94208, 56.73071, 56.76717, 57.12477, 57.8536, 58.94226, 
    60.28629, 61.69645, 62.9693, 64.08333, 64.80651, 65.17484,
  61.79995, 61.47795, 60.89214, 60.13709, 59.31602, 58.5196, 57.75945, 
    57.23611, 56.86794, 56.69021, 56.7615, 57.14008, 57.85917, 58.89492, 
    60.14524, 61.44362, 62.61606, 63.65982, 64.33743, 64.68681,
  61.11716, 60.8734, 60.40819, 59.76575, 59.01525, 58.24669, 57.4812, 
    56.95633, 56.60469, 56.4631, 56.57686, 56.98357, 57.6918, 58.65764, 
    59.77868, 60.91616, 61.93386, 62.85171, 63.43879, 63.74576,
  60.27107, 60.0988, 59.74297, 59.19969, 58.50362, 57.74159, 56.95282, 
    56.38852, 56.02086, 55.89411, 56.04173, 56.4798, 57.18783, 58.09451, 
    59.09003, 60.05909, 60.90112, 61.64207, 62.10386, 62.34728,
  59.37774, 59.25288, 58.96669, 58.47776, 57.79085, 56.98593, 56.14517, 
    55.46523, 55.01105, 54.84497, 54.99651, 55.46644, 56.20402, 57.09994, 
    58.02201, 58.86456, 59.55501, 60.08485, 60.41559, 60.58828,
  58.52, 58.42074, 58.16745, 57.68924, 56.96272, 56.05428, 55.12024, 
    54.20485, 53.55079, 53.25609, 53.36087, 53.86673, 54.69361, 55.67188, 
    56.61713, 57.41444, 58.01818, 58.33802, 58.5714, 58.6883,
  57.79332, 57.7002, 57.44674, 56.94067, 56.1353, 55.07725, 33.86139, 
    32.47908, 31.41851, 30.83251, 30.78826, 31.33193, 32.3716, 33.62815, 
    34.78964, 35.69132, 36.31931, 56.66047, 56.85428, 56.9447,
  57.19871, 57.11301, 56.8614, 56.32713, 55.43062, 54.18201, 32.48869, 
    30.47445, 28.80774, 27.73854, 27.42024, 28.00544, 29.39988, 31.13994, 
    32.70667, 33.87334, 34.68401, 55.20903, 55.44526, 55.55057,
  56.76562, 56.69349, 56.45554, 55.90963, 54.9417, 53.52279, 31.41047, 
    28.78606, 26.5149, 24.95305, 24.34554, 24.9603, 26.72853, 29.00603, 
    31.03609, 32.51163, 33.53381, 54.1772, 54.48013, 54.61679,
  56.53258, 56.48071, 56.27126, 55.7396, 54.74123, 53.21351, 30.80073, 
    27.68638, 24.91695, 22.96866, 22.15319, 22.79928, 24.87353, 27.61202, 
    30.04168, 31.77003, 32.9513, 53.67556, 54.03522, 54.20178,
  56.56291, 56.53262, 56.35791, 55.85902, 54.87199, 53.31526, 30.74434, 
    27.35219, 24.28771, 22.12956, 21.22347, 21.90533, 24.167, 27.19143, 
    29.86236, 31.72777, 32.98517, 53.77581, 54.17105, 54.35928,
  56.9258, 56.90887, 56.75846, 56.2915, 55.34169, 53.83078, 31.29633, 
    27.94802, 24.91437, 22.78959, 21.92061, 22.63894, 24.9311, 27.96675, 
    30.62125, 32.45706, 33.69228, 54.50924, 54.91828, 55.11928,
  57.66588, 57.64157, 57.48249, 57.01741, 56.09706, 54.66727, 32.36037, 
    29.37081, 26.71863, 24.90614, 24.22718, 24.97586, 27.09952, 29.82912, 
    32.20343, 33.86971, 35.01844, 55.80033, 56.21186, 56.42036,
  58.76569, 58.70198, 58.48033, 57.95756, 57.0182, 55.64336, 33.64474, 
    31.13877, 29.02801, 27.67747, 27.28257, 28.04164, 29.8611, 32.12947, 
    34.14156, 35.63433, 36.72148, 57.4326, 57.85327, 58.06973,
  60.12117, 59.98414, 59.641, 58.98966, 57.96023, 56.57339, 34.82654, 
    32.72806, 31.07891, 30.12043, 29.95959, 30.70175, 32.24481, 34.15157, 
    35.92944, 37.36229, 38.47182, 59.1254, 59.57162, 59.79985,
  61.55803, 61.32649, 60.82234, 59.98944, 58.80955, 57.34748, 35.73104, 
    33.9144, 32.57347, 31.85734, 31.82463, 32.53573, 33.91092, 35.64163, 
    37.35563, 38.83752, 40.02672, 60.65551, 61.13746, 61.38096,
  62.89228, 62.5658, 61.89401, 60.86089, 59.49993, 57.92687, 36.3274, 
    34.7308, 33.60632, 33.03802, 33.07079, 33.75555, 35.04334, 36.70963, 
    38.44237, 40.0031, 41.26282, 61.90014, 62.41904, 62.68148,
  63.97234, 63.57375, 62.76743, 61.56027, 60.02404, 58.32101, 56.7074, 
    55.28778, 54.28288, 53.7817, 53.85218, 54.54158, 55.80244, 57.43956, 
    59.16917, 60.7438, 62.00914, 62.78379, 63.35809, 63.65138,
  64.75063, 64.30354, 63.39947, 62.05587, 60.37717, 58.57123, 56.86427, 
    55.52003, 54.5817, 54.12263, 54.21683, 54.91839, 56.19082, 57.85163, 
    59.6164, 61.21983, 62.4933, 63.40973, 64.01459, 64.32743,
  65.18047, 64.7146, 63.76308, 62.33941, 60.56626, 58.68604, 56.91549, 
    55.59003, 54.6739, 54.22747, 54.32838, 55.04208, 56.34381, 58.05151, 
    59.86415, 61.49673, 62.77747, 63.75878, 64.3782, 64.70097,
  63.27683, 62.86745, 62.09785, 61.06108, 59.88324, 58.70237, 57.5879, 
    56.77346, 56.20602, 55.93409, 56.01934, 56.51132, 57.41646, 58.66522, 
    60.10517, 61.53769, 62.78744, 63.87326, 64.58042, 64.94582,
  62.82761, 62.46455, 61.77653, 60.83517, 59.74231, 58.62157, 57.53889, 
    56.74498, 56.19794, 55.95025, 56.05561, 56.5484, 57.41998, 58.59637, 
    59.93864, 61.27427, 62.44827, 63.48297, 64.15746, 64.50861,
  62.03734, 61.74833, 61.18835, 60.39409, 59.43096, 58.40143, 57.36641, 
    56.59444, 56.06825, 55.84906, 55.97978, 56.47276, 57.29666, 58.36891, 
    59.56681, 60.75313, 61.80233, 62.73759, 63.34561, 63.66554,
  60.98535, 60.78017, 60.36345, 59.73202, 58.91137, 57.97931, 57.00122, 
    56.23418, 55.71434, 55.51693, 55.6733, 56.16951, 56.94522, 57.90372, 
    58.93605, 59.9417, 60.82908, 61.60485, 62.11219, 62.38187,
  59.78862, 59.65775, 59.36706, 58.87734, 58.17713, 57.31774, 56.39458, 
    55.58208, 55.0249, 54.8214, 54.99431, 55.50238, 56.25006, 57.11704, 
    57.99928, 58.82693, 59.54297, 60.09823, 60.4841, 60.6898,
  58.57747, 58.50084, 58.30156, 57.91201, 57.28794, 56.45043, 55.5542, 
    54.5928, 53.9028, 53.62873, 53.79503, 54.33599, 55.1096, 55.95102, 
    56.74363, 57.43927, 58.01767, 58.32535, 58.60125, 58.74599,
  57.50969, 57.45959, 57.3047, 56.96122, 56.36121, 55.49144, 34.4287, 
    33.07704, 32.03083, 31.5319, 31.627, 32.24441, 33.17934, 34.16834, 
    35.03165, 35.72054, 36.2575, 56.531, 56.74208, 56.84698,
  56.64969, 56.61366, 56.48062, 56.15242, 55.53451, 54.5681, 33.0937, 
    31.17701, 29.54979, 28.60831, 28.50175, 29.21008, 30.44634, 31.76896, 
    32.87949, 33.72545, 34.38929, 54.91033, 55.15107, 55.26252,
  56.05952, 56.0336, 55.91564, 55.59557, 54.95559, 53.89368, 32.03827, 
    29.53985, 27.2682, 25.78759, 25.39564, 26.18598, 27.81113, 29.6019, 
    31.08505, 32.18565, 33.0483, 53.7636, 54.07189, 54.21286,
  55.78503, 55.77039, 55.67126, 55.36907, 54.72923, 53.61839, 31.52436, 
    28.57955, 25.76187, 23.80018, 23.14618, 24.01266, 26.01377, 28.25805, 
    30.08826, 31.40909, 32.43004, 53.26377, 53.63468, 53.80766,
  55.87822, 55.87247, 55.78988, 55.50895, 54.88872, 53.7846, 31.61623, 
    28.46814, 25.35759, 23.1298, 22.34295, 23.27614, 25.51826, 28.03544, 
    30.05339, 31.47692, 32.56559, 53.46232, 53.87239, 54.06965,
  56.38057, 56.37159, 56.28542, 56.00567, 55.39767, 54.32725, 32.24642, 
    29.18986, 26.1613, 24.01042, 23.2908, 24.26218, 26.49898, 28.97553, 
    30.9444, 32.33404, 33.40561, 54.29729, 54.72309, 54.93468,
  57.29094, 57.2557, 57.1254, 56.79821, 56.15795, 55.09613, 33.20107, 
    30.44335, 27.80756, 26.03529, 25.55544, 26.52058, 28.51561, 30.68605, 
    32.44233, 33.73532, 34.76498, 55.58736, 56.01771, 56.23654,
  58.53598, 58.44674, 58.22201, 57.78277, 57.0408, 55.92195, 34.20518, 
    31.77743, 29.61155, 28.28964, 28.0764, 28.99906, 30.68851, 32.51999, 
    34.08049, 35.32134, 36.34996, 57.07894, 57.51647, 57.73997,
  59.97026, 59.80638, 59.44767, 58.84119, 57.93257, 56.68933, 35.07134, 
    32.89724, 31.10671, 30.12541, 30.09186, 30.96264, 32.43736, 34.06895, 
    35.55413, 36.8221, 37.89698, 58.54628, 58.99768, 59.22641,
  61.41623, 61.17312, 60.66763, 59.86914, 58.75836, 57.35209, 35.74225, 
    33.75093, 32.22321, 31.45578, 31.51651, 32.34858, 33.72135, 35.29299, 
    36.80016, 38.13461, 39.26095, 59.85225, 60.31953, 60.55528,
  62.72011, 62.40756, 61.76774, 60.78348, 59.46733, 57.89099, 36.22577, 
    34.40562, 33.0917, 32.47619, 32.5949, 33.40345, 34.72934, 36.29466, 
    37.84465, 39.23054, 40.37413, 60.92866, 61.41014, 61.65603,
  63.76658, 63.40712, 62.66914, 61.53464, 60.03334, 58.2839, 56.5548, 
    54.93142, 53.78281, 53.26405, 53.42559, 54.22916, 55.52032, 57.05204, 
    58.58131, 59.94519, 61.05184, 61.69445, 62.21564, 62.4875,
  64.52175, 64.13366, 63.33009, 62.08627, 60.44419, 58.56345, 56.70398, 
    55.14834, 54.07704, 53.61529, 53.81245, 54.63614, 55.94231, 57.49109, 
    59.03457, 60.39863, 61.48747, 62.25269, 62.79613, 63.08508,
  64.93987, 64.54438, 63.71455, 62.41189, 60.67977, 58.70497, 56.75249, 
    55.20205, 54.15396, 53.71624, 53.93655, 54.78881, 56.13235, 57.71938, 
    59.28801, 60.65799, 61.73956, 62.56501, 63.12262, 63.42241,
  63.88606, 63.48082, 62.69034, 61.56627, 60.21106, 58.78099, 57.39919, 
    56.36061, 55.65992, 55.36316, 55.51539, 56.12218, 57.12976, 58.41571, 
    59.81088, 61.14406, 62.28576, 63.2884, 63.94898, 64.29661,
  63.43212, 63.05704, 62.32787, 61.29162, 60.03556, 58.69509, 57.37681, 
    56.375, 55.69503, 55.41003, 55.56134, 56.14424, 57.09793, 58.30568, 
    59.61636, 60.87803, 61.96878, 62.93374, 63.56838, 63.90305,
  62.61153, 62.29264, 61.67118, 60.78008, 59.68092, 58.47885, 57.26004, 
    56.30828, 55.65443, 55.38391, 55.53292, 56.0812, 56.95623, 58.04698, 
    59.22632, 60.37111, 61.37401, 62.26285, 62.84798, 63.15792,
  61.46978, 61.22706, 60.74624, 60.03714, 59.12896, 58.09217, 57.00269, 
    56.10038, 55.47087, 55.21616, 55.36551, 55.87796, 56.66342, 57.61362, 
    58.62716, 59.61558, 60.49357, 61.25059, 61.75992, 62.03122,
  60.10366, 59.94396, 59.613, 59.09288, 58.3785, 57.50404, 56.56202, 
    55.68051, 55.05285, 54.80507, 54.95897, 55.44686, 56.15233, 56.96281, 
    57.79961, 58.61, 59.33752, 59.89351, 60.30453, 60.52399,
  58.65922, 58.57381, 58.37585, 58.02145, 57.47272, 56.72535, 55.91629, 
    54.97535, 54.27656, 53.99624, 54.15541, 54.65006, 55.31845, 56.02778, 
    56.71478, 57.36075, 57.94447, 58.25177, 58.56104, 58.72441,
  57.33783, 57.30047, 57.19046, 56.94898, 56.51457, 55.84215, 34.97397, 
    33.74656, 32.7552, 32.30692, 32.44837, 33.02567, 33.78714, 34.53386, 
    35.19118, 35.76435, 36.27407, 56.51833, 56.7507, 56.86784,
  56.26882, 56.25723, 56.19482, 56.0132, 55.62972, 54.95435, 33.77048, 
    32.11902, 30.64579, 29.84112, 29.86059, 30.53531, 31.48848, 32.39949, 
    33.15281, 33.77817, 34.34818, 54.87313, 55.11655, 55.22994,
  55.56067, 55.55899, 55.51595, 55.3597, 54.99459, 54.29293, 32.78254, 
    30.65478, 28.58936, 27.27742, 27.06524, 27.84805, 29.11857, 30.36344, 
    31.36907, 32.17321, 32.90304, 53.68482, 53.98304, 54.11744,
  55.27364, 55.27365, 55.2359, 55.09019, 54.73653, 54.02572, 32.33224, 
    29.85195, 27.27609, 25.467, 24.99784, 25.88766, 27.51032, 29.12404, 
    30.39774, 31.38183, 32.25838, 53.18542, 53.54053, 53.70246,
  55.44051, 55.43355, 55.38612, 55.23466, 54.8843, 54.1854, 32.47924, 
    29.87909, 27.06696, 24.99623, 24.39221, 25.363, 27.20422, 29.02516, 
    30.43358, 31.50268, 32.44548, 53.41345, 53.80317, 53.98655,
  56.05636, 56.02779, 55.94402, 55.75306, 55.37335, 54.67143, 33.06977, 
    30.56341, 27.8555, 25.8878, 25.36203, 26.35306, 28.15702, 29.92332, 
    31.29806, 32.36296, 33.30866, 54.22635, 54.62806, 54.82324,
  57.06008, 56.99057, 56.83386, 56.55313, 56.08529, 55.32135, 33.84177, 
    31.51591, 29.12088, 27.50221, 27.19037, 28.14095, 29.73014, 31.29243, 
    32.56855, 33.61885, 34.56519, 55.37761, 55.78172, 55.98173,
  58.32985, 58.20307, 57.94053, 57.52077, 56.90129, 56.00256, 34.5867, 
    32.41676, 30.3553, 29.10435, 28.99481, 29.8848, 31.26418, 32.65571, 
    33.87806, 34.95386, 35.92914, 56.62773, 57.03514, 57.23731,
  59.70911, 59.51932, 59.1362, 58.54923, 57.73593, 56.65254, 35.22511, 
    33.15918, 31.35944, 30.37877, 30.39986, 31.24804, 32.5169, 33.84547, 
    35.08153, 36.2088, 37.22044, 57.8208, 58.23359, 58.43813,
  61.04879, 60.80193, 60.3049, 59.55091, 58.53433, 57.25262, 35.75616, 
    33.77189, 32.16973, 31.37241, 31.47376, 32.30883, 33.55011, 34.89138, 
    36.17228, 37.34104, 38.3638, 58.88252, 59.29932, 59.5075,
  62.238, 61.94543, 61.35296, 60.45107, 59.24667, 57.78034, 36.19048, 
    34.31068, 32.89463, 32.24739, 32.40958, 33.24027, 34.47374, 35.83563, 
    37.14743, 38.32605, 39.3216, 59.77303, 60.19004, 60.40339,
  63.19342, 62.87149, 62.21225, 61.19487, 59.82626, 58.18012, 56.49922, 
    54.811, 53.59045, 53.06252, 53.26535, 54.07629, 55.26308, 56.57852, 
    57.84581, 58.97136, 59.90084, 60.39707, 60.84237, 61.07768,
  63.88913, 63.54922, 62.84652, 61.74902, 60.26186, 58.48385, 56.65157, 
    55.01249, 53.86667, 53.40157, 53.64538, 54.47817, 55.6762, 56.9963, 
    58.2579, 59.36366, 60.25999, 60.86141, 61.32139, 61.57032,
  64.27787, 63.93384, 63.21547, 62.07808, 60.51875, 58.64824, 56.70589, 
    55.05375, 53.9229, 53.48701, 53.76685, 54.63902, 55.87362, 57.2177, 
    58.48542, 59.58307, 60.46472, 61.12114, 61.59242, 61.85064,
  63.94093, 63.5706, 62.83521, 61.75379, 60.38653, 58.86423, 57.32919, 
    56.1241, 55.31515, 55.00438, 55.21025, 55.86367, 56.831, 57.95383, 
    59.09082, 60.13697, 61.02209, 61.82383, 62.3578, 62.6451,
  63.51818, 63.16229, 62.46148, 61.44153, 60.16248, 58.74223, 57.30257, 
    56.16059, 55.38117, 55.06843, 55.24417, 55.84419, 56.74467, 57.80151, 
    58.88527, 59.89504, 60.75651, 61.53401, 62.05016, 62.32732,
  62.74764, 62.42339, 61.79077, 60.87996, 59.74592, 58.48536, 57.19536, 
    56.14466, 55.40824, 55.09408, 55.22813, 55.75191, 56.55352, 57.50768, 
    58.50338, 59.4498, 60.27055, 60.99839, 61.48428, 61.74458,
  61.65126, 61.37864, 60.85012, 60.0938, 59.15237, 58.0944, 57.00127, 
    56.05736, 55.37404, 55.06387, 55.15478, 55.59137, 56.27229, 57.09319, 
    57.96717, 58.82042, 59.57977, 60.21798, 60.66059, 60.89695,
  60.28978, 60.08698, 59.69303, 59.1253, 58.40635, 57.571, 56.7085, 55.86447, 
    55.23132, 54.93005, 54.98664, 55.34122, 55.89636, 56.56717, 57.29446, 
    58.02757, 58.70493, 59.19638, 59.58292, 59.7878,
  58.78221, 58.65828, 58.41227, 58.04415, 57.55043, 56.92723, 56.29272, 
    55.50209, 54.87812, 54.57222, 54.61018, 54.9109, 55.36264, 55.89286, 
    56.47132, 57.07477, 57.66253, 57.95742, 58.28053, 58.44833,
  57.32962, 57.27415, 57.15693, 56.96346, 56.66726, 56.22267, 35.63358, 
    34.72435, 33.93056, 33.52298, 33.55454, 33.88242, 34.32624, 34.79918, 
    35.29417, 35.8149, 36.34929, 56.61001, 56.87033, 56.9987,
  56.11494, 56.10554, 56.07545, 56.00054, 55.8368, 55.50249, 34.76088, 
    33.70887, 32.69443, 32.1125, 32.08501, 32.42168, 32.86293, 33.29505, 
    33.7253, 34.18651, 34.69902, 55.23841, 55.48849, 55.60357,
  55.31298, 55.32178, 55.32866, 55.30958, 55.21584, 54.94311, 33.99356, 
    32.73725, 31.41459, 30.55576, 30.41268, 30.78643, 31.3188, 31.82457, 
    32.29361, 32.78135, 33.34401, 54.17858, 54.44596, 54.56248,
  55.01619, 55.01915, 55.01923, 55.0004, 54.92041, 54.66956, 33.60642, 
    32.19469, 30.60518, 29.46458, 29.18272, 29.60291, 30.2713, 30.90633, 
    31.46879, 32.03278, 32.67775, 53.66319, 53.95605, 54.08203,
  55.22981, 55.20757, 55.16458, 55.09764, 54.97866, 54.70796, 33.65324, 
    32.18885, 30.48719, 29.20553, 28.84527, 29.29228, 30.04456, 30.7679, 
    31.4109, 32.05103, 32.7594, 53.73443, 54.042, 54.1768,
  55.87672, 55.81472, 55.69988, 55.54282, 55.33219, 54.98605, 33.9878, 
    32.51934, 30.84125, 29.5937, 29.2534, 29.69963, 30.45317, 31.20655, 
    31.91326, 32.62746, 33.38173, 54.24173, 54.55185, 54.69127,
  56.82328, 56.71375, 56.50944, 56.23149, 55.88298, 55.40112, 34.42228, 
    32.92787, 31.32261, 30.20293, 29.94217, 30.38281, 31.11042, 31.88197, 
    32.65734, 33.45235, 34.2528, 54.96797, 55.27721, 55.41865,
  57.91998, 57.76363, 57.46732, 57.05628, 56.54288, 55.88414, 34.86441, 
    33.31351, 31.77849, 30.79627, 30.62644, 31.08419, 31.8158, 32.6242, 
    33.46739, 34.33003, 35.16686, 55.7498, 56.05917, 56.20235,
  59.03949, 58.84364, 58.46609, 57.92937, 57.24959, 56.40496, 35.30672, 
    33.69586, 32.21635, 31.34698, 31.26275, 31.769, 32.54692, 33.40945, 
    34.30208, 35.19476, 36.03567, 56.50534, 56.81393, 56.95923,
  60.09136, 59.86555, 59.42366, 58.78115, 57.95364, 56.94062, 35.75206, 
    34.10641, 32.68422, 31.91319, 31.90994, 32.47791, 33.31603, 34.22818, 
    35.14171, 36.02243, 36.82775, 57.19843, 57.50182, 57.64878,
  61.01579, 60.76707, 60.2753, 59.54846, 58.60016, 57.44972, 36.18729, 
    34.5517, 33.21841, 32.55246, 32.61847, 33.22617, 34.09789, 35.03277, 
    35.94, 36.78089, 37.52082, 57.79907, 58.08944, 58.23591,
  61.75995, 61.49558, 60.96797, 60.17493, 59.12102, 57.83776, 56.50967, 
    55.0314, 53.89159, 53.34763, 53.43833, 54.00381, 54.81081, 55.6781, 
    56.5124, 57.27238, 57.9235, 58.18948, 58.4931, 58.65468,
  62.30812, 62.03257, 61.48055, 60.64359, 59.51934, 58.14464, 56.67999, 
    55.22418, 54.13451, 53.63939, 53.76221, 54.34054, 55.14624, 56.00077, 
    56.81072, 57.53639, 58.14405, 58.48864, 58.79503, 58.96356,
  62.61859, 62.33846, 61.77617, 60.91846, 59.75476, 58.31831, 56.75325, 
    55.26818, 54.17316, 53.6997, 53.86129, 54.47793, 55.30752, 56.1673, 
    56.96823, 57.67775, 58.26601, 58.65487, 58.96516, 59.13822,
  63.44963, 63.11478, 62.45416, 61.48516, 60.25108, 58.85184, 57.40467, 
    56.23513, 55.42893, 55.10437, 55.27084, 55.8319, 56.63599, 57.53609, 
    58.42508, 59.23406, 59.91562, 60.55087, 60.97271, 61.20252,
  63.0677, 62.74326, 62.10719, 61.18311, 60.01863, 58.70926, 57.3591, 
    56.26145, 55.49229, 55.16398, 55.29153, 55.79311, 56.5349, 57.38384, 
    58.23828, 59.02725, 59.69744, 60.3161, 60.72662, 60.94975,
  62.37686, 62.07446, 61.48679, 60.64404, 59.5965, 58.42947, 57.23199, 
    56.23847, 55.52422, 55.19364, 55.26836, 55.68546, 56.3346, 57.10271, 
    57.89886, 58.65319, 59.30616, 59.88982, 60.28217, 60.4944,
  61.39901, 61.13355, 60.62269, 59.90026, 59.01438, 58.03316, 57.03812, 
    56.16935, 55.52422, 55.19716, 55.21394, 55.53073, 56.06337, 56.72373, 
    57.43735, 58.14016, 58.76881, 59.28858, 59.65698, 59.85452,
  60.18097, 59.96926, 59.56518, 59.00002, 58.31195, 57.54413, 56.7887, 
    56.04749, 55.47618, 55.16, 55.12371, 55.33743, 55.74132, 56.27477, 
    56.88503, 57.51897, 58.11521, 58.52928, 58.86899, 59.04811,
  58.81304, 58.66887, 58.39451, 58.01116, 57.53879, 56.98811, 56.47461, 
    55.83617, 55.31827, 55.00958, 54.93203, 55.05728, 55.33994, 55.74519, 
    56.24479, 56.80074, 57.36123, 57.63342, 57.94101, 58.09807,
  57.46078, 57.38438, 57.23907, 57.03438, 56.77068, 56.4217, 35.98116, 
    35.3265, 34.7365, 34.36912, 34.26025, 34.34978, 34.56943, 34.89564, 
    35.32357, 35.83094, 36.38102, 56.67347, 56.94047, 57.069,
  56.29465, 56.2711, 56.22585, 56.15866, 56.05518, 55.86273, 35.37386, 
    34.76254, 34.15789, 33.75176, 33.58826, 33.59055, 33.69151, 33.8889, 
    34.19807, 34.61351, 35.11305, 55.65484, 55.90477, 56.01853,
  55.50084, 55.50277, 55.50763, 55.51436, 55.50648, 55.42031, 34.82535, 
    34.21941, 33.57656, 33.12189, 32.90916, 32.84556, 32.86372, 32.96998, 
    33.18793, 33.53024, 33.99459, 54.80832, 55.04624, 55.14827,
  55.18468, 55.18273, 55.18343, 55.19278, 55.20271, 55.15244, 34.49096, 
    33.87096, 33.19519, 32.70339, 32.45231, 32.33908, 32.30326, 32.36006, 
    32.53952, 32.86488, 33.33883, 54.28266, 54.51636, 54.61246,
  55.34474, 55.31527, 55.26674, 55.21625, 55.16946, 55.07621, 34.4005, 
    33.7336, 33.01491, 32.48419, 32.19675, 32.05194, 32.00553, 32.08278, 
    32.30996, 32.69538, 33.22006, 54.12906, 54.36202, 54.45677,
  55.88363, 55.81357, 55.68914, 55.53769, 55.37813, 55.17285, 34.48944, 
    33.71902, 32.91733, 32.3233, 31.99795, 31.85837, 31.87086, 32.05353, 
    32.4095, 32.91183, 33.50854, 54.28363, 54.51605, 54.61161,
  56.65761, 56.54516, 56.33859, 56.07077, 55.7693, 55.40855, 34.685, 
    33.76811, 32.86026, 32.20311, 31.86492, 31.77848, 31.89962, 32.22228, 
    32.72321, 33.34357, 34.00686, 54.62813, 54.86063, 54.95811,
  57.53125, 57.38264, 57.10334, 56.72591, 56.28066, 55.75368, 34.96177, 
    33.89646, 32.89139, 32.19571, 31.88481, 31.89213, 32.13892, 32.58432, 
    33.18808, 33.87974, 34.57737, 55.06201, 55.29446, 55.39452,
  58.40704, 58.23148, 57.89605, 57.42875, 56.85802, 56.18135, 35.31773, 
    34.13378, 33.05453, 32.34631, 32.0941, 32.21628, 32.58499, 33.11898, 
    33.76847, 34.47094, 35.15748, 55.52452, 55.75379, 55.85603,
  59.22333, 59.02889, 58.65341, 58.11917, 57.45053, 56.65538, 35.73351, 
    34.47507, 33.35595, 32.66233, 32.48239, 32.71082, 33.17576, 33.76134, 
    34.41127, 35.07837, 35.71406, 55.97788, 56.19765, 56.30008,
  59.93876, 59.72993, 59.32486, 58.74205, 58.00285, 57.12451, 36.17723, 
    34.88925, 33.7763, 33.12606, 33.01043, 33.3063, 33.82339, 34.42684, 
    35.05284, 35.66367, 36.22464, 56.38747, 56.58768, 56.68604,
  60.51223, 60.29264, 59.86494, 59.24229, 58.43929, 57.47898, 56.51794, 
    55.3601, 54.40742, 53.8561, 53.75263, 54.00076, 54.44807, 54.9752, 
    55.51795, 56.04014, 56.50628, 56.62333, 56.82725, 56.93578,
  60.93655, 60.70855, 60.26474, 59.61658, 58.77448, 57.7617, 56.69762, 
    55.55387, 54.62859, 54.10383, 54.01756, 54.2695, 54.70837, 55.21608, 
    55.72923, 56.21413, 56.63467, 56.81211, 57.01118, 57.12217,
  61.17841, 60.94571, 60.49356, 59.83277, 58.96933, 57.92106, 56.78082, 
    55.61206, 54.67178, 54.15472, 54.09496, 54.37402, 54.82682, 55.33323, 
    55.83468, 56.30263, 56.70245, 56.91589, 57.1137, 57.22601,
  62.06831, 61.80775, 61.30537, 60.58802, 59.69188, 58.67926, 57.60778, 
    56.71243, 56.03553, 55.67728, 55.65273, 55.89153, 56.28756, 56.74846, 
    57.21392, 57.64434, 58.00627, 58.37527, 58.61448, 58.74897,
  61.77848, 61.52572, 61.03935, 60.34822, 59.49216, 58.53536, 57.53523, 
    56.69995, 56.06208, 55.70773, 55.65437, 55.84869, 56.2031, 56.6354, 
    57.08632, 57.51282, 57.87709, 58.24061, 58.47876, 58.61235,
  61.26415, 61.02504, 60.56692, 59.92179, 59.13382, 58.26696, 57.3814, 
    56.63316, 56.05381, 55.70964, 55.61917, 55.75096, 56.04354, 56.43142, 
    56.85989, 57.28311, 57.65726, 58.00653, 58.24428, 58.37638,
  60.55386, 60.33572, 59.92076, 59.34439, 58.65404, 57.90922, 57.18008, 
    56.53991, 56.03554, 55.70813, 55.57413, 55.62701, 55.83854, 56.1668, 
    56.56559, 56.98717, 57.38129, 57.70304, 57.9436, 58.07449,
  59.68766, 59.50005, 59.14672, 58.66496, 58.10193, 57.50658, 56.96951, 
    56.45266, 56.03747, 55.73489, 55.55374, 55.51348, 55.62593, 55.87989, 
    56.24148, 56.66193, 57.08593, 57.36345, 57.61185, 57.74207,
  58.72226, 58.57611, 58.30431, 57.94225, 57.53137, 57.10375, 56.76988, 
    56.38699, 56.07321, 55.80374, 55.57216, 55.42499, 55.42276, 55.59167, 
    55.9113, 56.33068, 56.7911, 57.01628, 57.27387, 57.40188,
  57.7536, 57.6557, 57.47757, 57.25033, 57.0069, 56.75869, 36.49646, 
    36.22331, 35.98738, 35.73867, 35.4456, 35.17646, 35.04873, 35.13334, 
    35.42276, 35.85768, 36.37169, 56.70203, 56.94905, 57.06348,
  56.87402, 56.82122, 56.72929, 56.62435, 56.53459, 56.4656, 36.28995, 
    36.28572, 36.30558, 36.20443, 35.86932, 35.39859, 35.02383, 34.9005, 
    35.04115, 35.37562, 35.82082, 56.31845, 56.53958, 56.63811,
  56.21096, 56.18783, 56.15284, 56.13087, 56.15282, 56.23147, 36.11234, 
    36.3809, 36.70573, 36.83364, 36.52327, 35.86974, 35.22313, 34.83855, 
    34.76, 34.91867, 35.22536, 55.89592, 56.06614, 56.1376,
  55.84687, 55.83035, 55.80818, 55.80725, 55.8652, 56.00597, 35.9053, 
    36.34256, 36.90876, 37.25354, 36.9961, 36.20193, 35.31907, 34.70085, 
    34.4305, 34.44392, 34.647, 55.39421, 55.52119, 55.5685,
  55.79263, 55.76146, 55.71068, 55.67006, 55.68289, 55.77778, 35.62953, 
    36.03268, 36.62863, 37.0261, 36.7652, 35.8901, 34.90437, 34.21568, 
    33.91734, 33.92845, 34.14038, 54.85581, 54.9673, 55.00291,
  55.98998, 55.93275, 55.83039, 55.71395, 55.62824, 55.59908, 35.34906, 
    35.53791, 35.93694, 36.18385, 35.83907, 34.96028, 34.05104, 33.49443, 
    33.34367, 33.48186, 33.78571, 54.39465, 54.51051, 54.54549,
  56.34897, 56.26503, 56.10921, 55.91151, 55.71428, 55.53869, 35.1783, 
    35.0941, 35.19865, 35.2005, 34.75401, 33.95187, 33.23649, 32.90219, 
    32.94618, 33.22805, 33.62398, 54.09821, 54.22163, 54.26064,
  56.78667, 56.68166, 56.48366, 56.22033, 55.92942, 55.62964, 35.19084, 
    34.87627, 34.70915, 34.48418, 33.97714, 33.306, 32.8058, 32.66259, 
    32.83843, 33.1991, 33.6363, 53.97792, 54.10291, 54.14567,
  57.2439, 57.12478, 56.89935, 56.59334, 56.23982, 55.85722, 35.38734, 
    34.91709, 34.54213, 34.14899, 33.63021, 33.10366, 32.78326, 32.76029, 
    32.98542, 33.35089, 33.7733, 53.99421, 54.11247, 54.15631,
  57.68064, 57.55299, 57.3125, 56.98469, 56.59945, 56.17579, 35.71679, 
    35.1536, 34.63225, 34.12815, 33.6263, 33.22382, 33.02971, 33.06704, 
    33.28653, 33.61001, 33.97862, 54.09363, 54.19638, 54.23736,
  58.06659, 57.93332, 57.685, 57.34981, 56.95793, 56.52977, 36.12487, 
    35.50322, 34.88083, 34.31169, 33.83796, 33.5256, 33.40934, 33.47074, 
    33.66231, 33.9268, 34.22139, 54.22767, 54.30307, 54.33517,
  58.37072, 58.23264, 57.97717, 57.63391, 57.23359, 56.80097, 56.4712, 
    55.93448, 55.39226, 54.86358, 54.39109, 54.04691, 53.87304, 53.85866, 
    53.96308, 54.13726, 54.33497, 54.25122, 54.31645, 54.35144,
  58.59848, 58.45645, 58.19592, 57.84943, 57.4491, 57.01904, 56.64312, 
    56.11632, 55.56913, 55.02909, 54.54984, 54.2006, 54.01535, 53.97944, 
    54.05303, 54.19012, 54.34248, 54.29157, 54.34196, 54.37363,
  58.72949, 58.58433, 58.3195, 57.96982, 57.56801, 57.1359, 56.72522, 
    56.19388, 55.63031, 55.07486, 54.59165, 54.24615, 54.06327, 54.02351, 
    54.0867, 54.20825, 54.33952, 54.31232, 54.35526, 54.38458,
  60.83565, 60.63912, 60.26886, 59.75722, 59.14038, 58.46355, 57.74481, 
    57.13721, 56.61582, 56.23751, 56.02748, 55.97052, 56.02773, 56.1576, 
    56.32595, 56.50205, 56.65455, 56.85073, 56.97249, 57.04587,
  60.62548, 60.43491, 60.07587, 59.58058, 58.98658, 58.34079, 57.66595, 
    57.09644, 56.6061, 56.23945, 56.01923, 55.9395, 55.97387, 56.08877, 
    56.25206, 56.43177, 56.59389, 56.79137, 56.91814, 56.99398,
  60.25977, 60.07826, 59.73674, 59.26797, 58.71177, 58.11616, 57.5146, 
    57.00152, 56.55959, 56.21468, 55.98355, 55.87213, 55.87291, 55.96632, 
    56.12537, 56.31709, 56.50342, 56.69984, 56.83702, 56.91714,
  59.76953, 59.60062, 59.28399, 58.8537, 58.35233, 57.82724, 57.33052, 
    56.89208, 56.51545, 56.20087, 55.9552, 55.7996, 55.75337, 55.81793, 
    55.97441, 56.18854, 56.41715, 56.60902, 56.76476, 56.85173,
  59.19249, 59.04092, 58.75884, 58.38204, 57.95547, 57.52305, 57.16247, 
    56.82158, 56.53152, 56.2576, 55.99098, 55.7725, 55.65952, 55.68364, 
    55.83675, 56.0817, 56.36948, 56.55563, 56.73875, 56.83469,
  58.56847, 58.4406, 58.20536, 57.89959, 57.56919, 57.25252, 57.04577, 
    56.83702, 56.66754, 56.45161, 56.15383, 55.84238, 55.63242, 55.59867, 
    55.74411, 56.02316, 56.37807, 56.56671, 56.77755, 56.88033,
  57.94833, 57.85009, 57.67326, 57.45541, 57.24288, 57.06792, 36.91895, 
    36.88051, 36.87225, 36.73742, 36.38995, 35.93229, 35.57103, 35.44923, 
    35.58273, 35.90466, 36.33543, 56.66138, 56.87075, 56.96488,
  57.35505, 57.28797, 57.17171, 57.04441, 56.95731, 56.95237, 36.95983, 
    37.28325, 37.6388, 37.73307, 37.37854, 36.70922, 36.06834, 35.71352, 
    35.69078, 35.91059, 36.26051, 56.67706, 56.85066, 56.92585,
  56.84231, 56.80131, 56.73531, 56.68326, 56.70414, 56.858, 37.01531, 
    37.71414, 38.4753, 38.86271, 38.56476, 37.7163, 36.77674, 36.12238, 
    35.84766, 35.8604, 36.0314, 56.53312, 56.63728, 56.67876,
  56.44998, 56.4231, 56.38305, 56.36816, 56.44279, 56.68153, 36.91993, 
    37.86216, 38.92421, 39.5503, 39.31626, 38.33925, 37.15287, 36.22862, 
    35.7145, 35.53049, 35.54635, 56.08617, 56.13214, 56.14376,
  56.20239, 56.17537, 56.13258, 56.10958, 56.16967, 56.38736, 36.58488, 
    37.52695, 38.64861, 39.33808, 39.10257, 38.04107, 36.72481, 35.67806, 
    35.074, 34.83161, 34.82041, 55.35144, 55.37988, 55.3782,
  56.09974, 56.06229, 55.99665, 55.93386, 55.92998, 56.04606, 36.11029, 
    36.83351, 37.7658, 38.31995, 37.99891, 36.89906, 35.60114, 34.6249, 
    34.11628, 33.96726, 34.04286, 54.51731, 54.55881, 54.5587,
  56.11951, 56.06823, 55.97393, 55.86308, 55.78195, 55.77488, 35.69786, 
    36.12112, 36.73622, 37.03697, 36.58919, 35.51063, 34.35368, 33.56982, 
    33.24276, 33.23644, 33.41856, 53.79556, 53.85399, 53.86081,
  56.22689, 56.16378, 56.04633, 55.89811, 55.75672, 55.65429, 35.49397, 
    35.66294, 35.96677, 36.00113, 35.44107, 34.43825, 33.47246, 32.88606, 
    32.7059, 32.79324, 33.03212, 53.29073, 53.35447, 53.36617,
  56.38582, 56.3152, 56.18494, 56.01817, 55.84682, 55.6963, 35.5261, 35.5293, 
    35.58739, 35.39968, 34.76555, 33.86285, 33.07225, 32.62497, 32.51465, 
    32.62267, 32.85752, 52.99668, 53.05239, 53.06425,
  56.56356, 56.48975, 56.35674, 56.18979, 56.01841, 55.86428, 35.7395, 
    35.64469, 35.51968, 35.16376, 34.48971, 33.68279, 33.0239, 32.65555, 
    32.55693, 32.63607, 32.82515, 52.85719, 52.89392, 52.90086,
  56.73155, 56.65729, 56.52815, 56.37438, 56.2273, 56.10634, 36.07046, 
    35.90331, 35.6306, 35.15233, 34.46864, 33.7485, 33.18461, 32.85827, 
    32.74451, 32.77388, 32.89516, 52.8138, 52.81897, 52.81438,
  56.86121, 56.78626, 56.65944, 56.51535, 56.38994, 56.30678, 56.38985, 
    56.26926, 56.01748, 55.53896, 54.85476, 54.12699, 53.52925, 53.13945, 
    52.94332, 52.88537, 52.9104, 52.7121, 52.69777, 52.6913,
  56.96331, 56.88782, 56.76328, 56.62877, 56.52384, 56.47117, 56.53645, 
    56.42006, 56.14555, 55.63659, 54.93535, 54.20266, 53.59784, 53.18998, 
    52.96508, 52.87175, 52.85272, 52.66843, 52.63341, 52.6204,
  57.02315, 56.94634, 56.82108, 56.68927, 56.59287, 56.55426, 56.60619, 
    56.49734, 56.21048, 55.67669, 54.95392, 54.21083, 53.60278, 53.1913, 
    52.95803, 52.85085, 52.8115, 52.64311, 52.59768, 52.58067,
  59.46766, 59.34415, 59.12122, 58.8329, 58.51312, 58.191, 57.84788, 
    57.55557, 57.21608, 56.83224, 56.43525, 56.07062, 55.77592, 55.56665, 
    55.4366, 55.36345, 55.31662, 55.35229, 55.3674, 55.3859,
  59.34754, 59.22748, 59.0104, 58.72908, 58.41681, 58.10289, 57.77542, 
    57.49551, 57.17418, 56.80798, 56.42161, 56.0591, 55.76178, 55.5507, 
    55.42388, 55.36061, 55.32949, 55.37246, 55.39758, 55.42126,
  59.14652, 59.03065, 58.82068, 58.54828, 58.24697, 57.94668, 57.65053, 
    57.39248, 57.10373, 56.76834, 56.39941, 56.0395, 55.73791, 55.52641, 
    55.41023, 55.37096, 55.37554, 55.42958, 55.47434, 55.50712,
  58.89502, 58.78392, 58.58229, 58.32162, 58.03701, 57.75929, 57.51497, 
    57.29376, 57.05515, 56.7626, 56.41251, 56.04827, 55.73457, 55.52074, 
    55.42212, 55.42216, 55.48508, 55.55533, 55.63138, 55.67749,
  58.625, 58.51964, 58.32881, 58.08523, 57.82763, 57.58836, 57.42124, 
    57.26601, 57.10604, 56.87167, 56.53589, 56.14817, 55.8017, 55.57419, 
    55.49406, 55.54404, 55.6835, 55.78144, 55.89833, 55.96012,
  58.35778, 58.26047, 58.08549, 57.86846, 57.65393, 57.4784, 57.41113, 
    57.37602, 57.34615, 57.19723, 56.86626, 56.41763, 55.9973, 55.72987, 
    55.65904, 55.75903, 55.97756, 56.12149, 56.27478, 56.34789,
  58.10163, 58.01632, 57.86589, 57.69049, 57.54275, 57.46659, 37.44228, 
    37.61289, 37.79677, 37.78107, 37.44074, 36.86404, 36.29008, 35.92784, 
    35.84511, 35.99186, 36.28459, 56.56683, 56.71738, 56.78189,
  57.81315, 57.7439, 57.62613, 57.50587, 57.44942, 57.52311, 37.70257, 
    38.26542, 38.83875, 39.07878, 38.77931, 38.04614, 37.22347, 36.63335, 
    36.38999, 36.42522, 36.61875, 56.9061, 57.00859, 57.04946,
  57.47184, 57.42213, 57.34296, 57.28457, 57.32602, 57.5587, 37.95109, 
    38.91008, 39.87327, 40.37733, 40.14945, 39.29944, 38.23656, 37.37428, 
    36.88461, 36.70594, 36.70321, 56.99083, 57.01305, 57.01652,
  57.06943, 57.0386, 56.99464, 56.98689, 57.09969, 57.44025, 37.968, 
    39.19152, 40.42406, 41.111, 40.93404, 40.00021, 38.74483, 37.63786, 
    36.90599, 36.51325, 36.33249, 56.62424, 56.58283, 56.55542,
  56.63704, 56.61944, 56.59793, 56.61581, 56.75205, 57.1111, 37.63246, 
    38.90262, 40.2089, 40.94632, 40.76028, 39.74751, 38.35563, 37.09119, 
    36.21773, 35.71825, 35.47839, 55.78689, 55.72996, 55.69106,
  56.23149, 56.2192, 56.20458, 56.22232, 56.33793, 56.63625, 37.03378, 
    38.14485, 39.32718, 39.97647, 39.71152, 38.61644, 37.15659, 35.86209, 
    34.99817, 34.53661, 34.364, 54.67629, 54.64254, 54.60928,
  55.90219, 55.88914, 55.87094, 55.8746, 55.94989, 56.15635, 36.40412, 
    37.25305, 38.18187, 38.63544, 38.23833, 37.07872, 35.63935, 34.43996, 
    33.70272, 33.36432, 33.30654, 53.57763, 53.57358, 53.5517,
  55.66918, 55.65337, 55.62986, 55.62111, 55.66409, 55.79782, 35.95428, 
    36.55809, 37.20468, 37.41647, 36.8714, 35.68867, 34.34654, 33.30387, 
    32.71446, 32.48726, 32.50924, 52.69228, 52.70168, 52.68723,
  55.52462, 55.50758, 55.48387, 55.47509, 55.51031, 55.61563, 35.76615, 
    36.19994, 36.60304, 36.58414, 35.91004, 34.74459, 33.52979, 32.6317, 
    32.1418, 31.96452, 32.00378, 52.07615, 52.07926, 52.06507,
  55.44511, 55.43, 55.4139, 55.42065, 55.47591, 55.59755, 35.80574, 36.13111, 
    36.33818, 36.12507, 35.35769, 34.23512, 33.13946, 32.34358, 31.89716, 
    31.71613, 31.72469, 51.68993, 51.67203, 51.6514,
  55.40324, 55.3927, 55.3907, 55.42626, 55.52611, 55.70145, 36.00852, 
    36.24321, 36.27675, 35.90792, 35.09349, 34.03944, 33.05155, 32.32507, 
    31.88805, 31.67397, 31.62422, 51.47055, 51.41743, 51.38307,
  55.3696, 55.36265, 55.37201, 55.4325, 55.57746, 55.81986, 56.26692, 
    56.50277, 56.50428, 56.10239, 55.28688, 54.25236, 53.26514, 52.49954, 
    51.99239, 51.69679, 51.55173, 51.25448, 51.17201, 51.13092,
  55.3565, 55.35258, 55.37147, 55.45284, 55.6341, 55.92538, 56.37043, 
    56.59876, 56.56311, 56.11988, 55.2835, 54.24894, 53.26395, 52.4882, 
    51.95702, 51.62884, 51.44128, 51.13803, 51.02916, 50.9785,
  55.35056, 55.34741, 55.3696, 55.45971, 55.65812, 55.97508, 56.42041, 
    56.66152, 56.61694, 56.14653, 55.27979, 54.22531, 53.23226, 52.4527, 
    51.91486, 51.57467, 51.36808, 51.07302, 50.95135, 50.89544,
  58.06578, 58.02053, 57.95299, 57.89431, 57.87038, 57.88992, 57.89891, 
    57.90004, 57.73846, 57.37041, 56.82387, 56.18714, 55.56327, 55.02588, 
    54.60403, 54.28999, 54.0562, 53.94637, 53.86768, 53.83875,
  58.04076, 57.99598, 57.92835, 57.86736, 57.83718, 57.8457, 57.84671, 
    57.83837, 57.68222, 57.33432, 56.81473, 56.20205, 55.59464, 55.06834, 
    54.65752, 54.35863, 54.14516, 54.04737, 53.98237, 53.96051,
  58.01197, 57.96613, 57.89504, 57.82656, 57.78422, 57.77641, 57.77407, 
    57.75929, 57.62074, 57.30836, 56.82839, 56.24779, 55.66248, 55.15444, 
    54.76651, 54.50052, 54.33088, 54.25444, 54.21601, 54.2068,
  58.00457, 57.9559, 57.87785, 57.79771, 57.74039, 57.71656, 57.7222, 
    57.71378, 57.61166, 57.35116, 56.91828, 56.36867, 55.80174, 55.31236, 
    54.95538, 54.73831, 54.63572, 54.59225, 54.59337, 54.60164,
  58.03859, 57.98555, 57.89812, 57.80512, 57.73624, 57.70747, 57.73986, 
    57.7706, 57.7386, 57.55151, 57.16754, 56.63403, 56.06543, 55.58093, 
    55.25221, 55.09077, 55.06867, 55.07774, 55.12528, 55.15207,
  58.11131, 58.05386, 57.95784, 57.85635, 57.7883, 57.78073, 57.864, 
    57.99789, 58.09491, 58.01522, 57.6784, 57.12876, 56.51542, 56.00162, 
    55.68233, 55.56686, 55.61638, 55.69838, 55.78075, 55.81857,
  58.19016, 58.13131, 58.03394, 57.93808, 57.89518, 57.94894, 38.06326, 
    38.4076, 38.729, 38.81077, 38.51843, 37.89946, 37.16503, 36.55718, 
    36.2109, 36.12241, 36.2218, 56.41297, 56.48404, 56.50989,
  58.17863, 58.12421, 58.03787, 57.96917, 57.98814, 58.1666, 38.50377, 
    39.20368, 39.86232, 40.17419, 39.96572, 39.28772, 38.39589, 37.60513, 
    37.10313, 36.88822, 36.86663, 56.98012, 56.9919, 56.98938,
  58.00177, 57.96057, 57.90191, 57.88255, 57.98805, 58.31551, 38.88757, 
    39.92874, 40.88408, 41.3841, 41.24868, 40.53624, 39.51245, 38.52796, 
    37.8171, 37.4002, 37.18373, 57.22777, 57.15611, 57.11528,
  57.61385, 57.59294, 57.57348, 57.61308, 57.80318, 58.25465, 38.99367, 
    40.2716, 41.42001, 42.02829, 41.92405, 41.17324, 40.0333, 38.86631, 
    37.9453, 37.32573, 36.93297, 56.95359, 56.81963, 56.74984,
  57.04211, 57.04307, 57.0636, 57.15523, 57.40339, 57.9158, 38.69735, 
    40.06474, 41.28881, 41.92823, 41.80381, 40.97921, 39.70869, 38.37269, 
    37.28279, 36.52793, 36.0542, 56.10863, 55.96199, 55.88382,
  56.37712, 56.39561, 56.44678, 56.57201, 56.84148, 57.34408, 38.05081, 
    39.35944, 40.54454, 41.1431, 40.94527, 40.00188, 38.58601, 37.1199, 
    35.9484, 35.17013, 34.73438, 54.84718, 54.73193, 54.66397,
  55.72534, 55.75458, 55.824, 55.96481, 56.2285, 56.67724, 37.25832, 
    38.40242, 39.44763, 39.92996, 39.60598, 38.51963, 36.98734, 35.47906, 
    34.34182, 33.64505, 33.32107, 53.46085, 53.3898, 53.33905,
  55.16264, 55.19781, 55.27795, 55.42702, 55.68007, 56.07433, 36.56173, 
    37.51182, 38.35793, 38.66245, 38.17739, 36.96541, 35.39273, 33.94385, 
    32.92068, 32.34182, 32.12273, 52.22561, 52.18191, 52.14352,
  54.7187, 54.7588, 54.84975, 55.0122, 55.26974, 55.64135, 36.11065, 
    36.89834, 37.53815, 37.64095, 36.99496, 35.70647, 34.17086, 32.83626, 
    31.93244, 31.43797, 31.26721, 51.2827, 51.23997, 51.2041,
  54.38748, 54.43436, 54.54151, 54.72967, 55.01587, 55.40587, 35.92051, 
    36.5849, 37.03499, 36.94682, 36.17213, 34.86352, 33.40991, 32.19022, 
    31.36748, 30.90403, 30.72551, 50.63854, 50.57566, 50.53312,
  54.14563, 54.20177, 54.33144, 54.55868, 54.89844, 55.34432, 35.94262, 
    36.49371, 36.76208, 36.50858, 35.65823, 34.38892, 33.04461, 31.92455, 
    31.14578, 30.67382, 30.45034, 50.23846, 50.13754, 50.07956,
  53.96119, 54.0251, 54.17432, 54.43853, 54.83877, 55.3654, 56.10129, 
    56.60552, 56.80042, 56.49129, 55.63754, 54.40987, 53.10598, 51.9842, 
    51.15818, 50.61494, 50.29756, 49.91405, 49.77285, 49.70298,
  53.84417, 53.91462, 54.08006, 54.37444, 54.82135, 55.40498, 56.14378, 
    56.6246, 56.77168, 56.41737, 55.54359, 54.323, 53.03417, 51.91506, 
    51.07352, 50.50207, 50.14377, 49.73208, 49.55836, 49.47583,
  53.7793, 53.85261, 54.02543, 54.33432, 54.80539, 55.4218, 56.16699, 
    56.65818, 56.79677, 56.41806, 55.51459, 54.27126, 52.97133, 51.84784, 
    51.00109, 50.4197, 50.04403, 49.63233, 49.44367, 49.35481,
  56.10427, 56.17767, 56.34139, 56.61256, 56.99058, 57.4415, 57.86281, 
    58.19149, 58.24163, 57.93592, 57.28308, 56.37994, 55.3753, 54.41281, 
    53.58728, 52.9331, 52.43998, 52.13662, 51.93805, 51.85009,
  56.22071, 56.2898, 56.44413, 56.69945, 57.05399, 57.47412, 57.86686, 
    58.17024, 58.21568, 57.92883, 57.31247, 56.45159, 55.48412, 54.54964, 
    53.74588, 53.11261, 52.64322, 52.35592, 52.17342, 52.09361,
  56.44404, 56.50426, 56.64011, 56.86684, 57.18354, 57.55953, 57.92016, 
    58.19847, 58.25083, 58.00051, 57.43816, 56.63362, 55.71428, 54.81843, 
    54.0498, 53.45563, 53.03371, 52.77698, 52.62514, 52.55984,
  56.78167, 56.82895, 56.93863, 57.12697, 57.39681, 57.72324, 58.05444, 
    58.31934, 58.39847, 58.20582, 57.71329, 56.97266, 56.10278, 55.24566, 
    54.51583, 53.9703, 53.61179, 53.40104, 53.28966, 53.24215,
  57.22135, 57.25316, 57.33228, 57.47834, 57.70154, 57.98652, 58.29629, 
    58.57792, 58.71514, 58.60528, 58.19612, 57.51911, 56.68736, 55.85353, 
    55.14983, 54.64562, 54.34775, 54.20419, 54.13112, 54.09851,
  57.71406, 57.7307, 57.78064, 57.88935, 58.07811, 58.34685, 58.65271, 
    59.00558, 59.24558, 59.24745, 58.93334, 58.31321, 57.49621, 56.65361, 
    55.94444, 55.4526, 55.18549, 55.11973, 55.06429, 55.03561,
  58.17542, 58.1816, 58.21246, 58.30066, 58.47948, 58.76765, 39.09154, 
    39.6045, 40.00988, 40.15649, 39.94833, 39.37729, 38.54679, 37.65322, 
    36.89669, 36.37882, 36.10018, 56.0652, 55.98335, 55.93641,
  58.46674, 58.4707, 58.50003, 58.59709, 58.81071, 59.18066, 39.70151, 
    40.42482, 41.01077, 41.29894, 41.20628, 40.71713, 39.906, 38.95607, 
    38.08869, 37.43488, 37.01204, 56.8019, 56.65277, 56.57381,
  58.48357, 58.4964, 58.54601, 58.68251, 58.96594, 59.44875, 40.16359, 
    41.07096, 41.78397, 42.15104, 42.12367, 41.6937, 40.90503, 39.90871, 
    38.92695, 38.11747, 37.52662, 57.17989, 56.95365, 56.83918,
  58.15834, 58.19004, 58.27831, 58.47652, 58.84893, 59.45225, 40.32539, 
    41.38195, 42.17934, 42.57698, 42.56043, 42.13376, 41.32038, 40.24683, 
    39.13733, 38.17627, 37.4391, 57.0386, 56.75783, 56.61901,
  57.49934, 57.55597, 57.69281, 57.96099, 58.42166, 59.12892, 40.10304, 
    41.28236, 42.14913, 42.55815, 42.50957, 42.01449, 41.09172, 39.87131, 
    38.60255, 37.50399, 36.67395, 56.30807, 56.01567, 55.87182,
  56.59404, 56.67601, 56.86039, 57.19117, 57.71977, 58.49133, 39.49625, 
    40.76088, 41.68605, 42.0976, 41.98073, 41.34404, 40.2224, 38.78786, 
    37.34489, 36.14947, 35.30811, 55.04551, 54.78747, 54.65814,
  55.58013, 55.6832, 55.90585, 56.28202, 56.84846, 57.63474, 38.60585, 
    39.8902, 40.83707, 41.2266, 41.00318, 40.16753, 38.79618, 37.13934, 
    35.56949, 34.35911, 33.59517, 53.45344, 53.25697, 53.15351,
  54.59591, 54.71467, 54.96516, 55.37105, 55.9523, 56.71854, 37.62823, 
    38.8554, 39.75937, 40.07962, 39.71405, 38.66243, 37.06595, 35.26488, 
    33.67389, 32.53719, 31.89744, 51.82718, 51.68673, 51.60727,
  53.73814, 53.86937, 54.14252, 54.5728, 55.16451, 55.90709, 36.77605, 
    37.89258, 38.68904, 38.89022, 38.36777, 37.13768, 35.41076, 33.58833, 
    32.07278, 31.04626, 30.50889, 50.42718, 50.31246, 50.24495,
  53.04796, 53.19168, 53.48904, 53.94948, 54.56457, 55.30523, 36.17095, 
    37.1548, 37.80281, 37.8577, 37.19626, 35.86445, 34.12045, 32.37225, 
    30.96702, 30.02737, 29.53298, 49.37902, 49.25572, 49.18563,
  52.52273, 52.68093, 53.0081, 53.51104, 54.17185, 54.9424, 35.83595, 
    36.67836, 37.1586, 37.06572, 36.30855, 34.96391, 33.29778, 31.67396, 
    30.37057, 29.47448, 28.96752, 48.68579, 48.52403, 48.43773,
  52.13046, 52.30157, 52.657, 53.20604, 53.93187, 54.77388, 55.77129, 
    56.50436, 56.87355, 56.7074, 55.93738, 54.64544, 53.06842, 51.51453, 
    50.22383, 49.28834, 48.69514, 48.19563, 47.97497, 47.86812,
  51.87473, 52.05676, 52.43584, 53.02252, 53.79787, 54.69056, 55.68913, 
    56.37523, 56.68755, 56.47753, 55.69106, 54.41473, 52.87273, 51.34883, 
    50.06573, 49.11492, 48.48459, 47.91754, 47.65371, 47.52901,
  51.73232, 51.92011, 52.312, 52.92006, 53.72552, 54.65302, 55.65804, 
    56.3428, 56.64301, 56.41557, 55.61033, 54.318, 52.76628, 51.23849, 
    49.95259, 48.99527, 48.35012, 47.76849, 47.48616, 47.35348,
  55.01988, 55.16701, 55.47067, 55.93145, 56.52234, 57.17714, 57.77089, 
    58.226, 58.36852, 58.12152, 57.47837, 56.51249, 55.36385, 54.19648, 
    53.146, 52.2867, 51.63283, 51.21152, 50.9415, 50.81914,
  55.22241, 55.36219, 55.6507, 56.08801, 56.64756, 57.26573, 57.82784, 
    58.25865, 58.39689, 58.16698, 57.55822, 56.63583, 55.53006, 54.3981, 
    53.37483, 52.53844, 51.90775, 51.50261, 51.24762, 51.13264,
  55.59432, 55.72094, 55.98325, 56.38246, 56.89538, 57.46383, 57.99029, 
    58.39859, 58.54482, 58.35026, 57.79467, 56.93134, 55.88011, 54.7933, 
    53.80803, 53.00895, 52.42097, 52.0466, 51.81939, 51.71717,
  56.12387, 56.2331, 56.46132, 56.8128, 57.27049, 57.7843, 58.27445, 
    58.67064, 58.84224, 58.70342, 58.21971, 57.42846, 56.43765, 55.39659, 
    54.44878, 53.68896, 53.15026, 52.82002, 52.62514, 52.53654,
  56.77036, 56.86078, 57.05265, 57.35495, 57.75914, 58.22575, 58.67928, 
    59.0851, 59.30334, 59.24008, 58.84542, 58.13704, 57.20708, 56.20178, 
    55.27555, 54.53831, 54.03372, 53.76413, 53.59288, 53.51244,
  57.45387, 57.52793, 57.6885, 57.95017, 58.31424, 58.75513, 59.18033, 
    59.6314, 59.92, 59.94875, 59.65746, 59.04172, 58.17017, 57.1821, 
    56.24699, 55.49593, 54.98612, 54.77768, 54.60842, 54.52544,
  58.06974, 58.1342, 58.27662, 58.51638, 58.86201, 59.30235, 39.7384, 
    40.29282, 40.68186, 40.81599, 40.64031, 40.13148, 39.32347, 38.33862, 
    37.36438, 36.55949, 35.99863, 55.76656, 55.56646, 55.46347,
  58.477, 58.54107, 58.68453, 58.9327, 59.30205, 59.79227, 40.38459, 
    41.04012, 41.50882, 41.72636, 41.66389, 41.2879, 40.5855, 39.63073, 
    38.59903, 37.6747, 36.97063, 56.52437, 56.25939, 56.1253,
  58.57928, 58.65299, 58.81734, 59.10196, 59.52681, 60.09375, 40.82623, 
    41.56537, 42.07886, 42.33146, 42.32848, 42.03969, 41.41845, 40.49272, 
    39.41395, 38.37889, 37.53619, 56.9317, 56.59837, 56.4324,
  58.31248, 58.40395, 58.60497, 58.94732, 59.45112, 60.11582, 40.97323, 
    41.80449, 42.35855, 42.62017, 42.6246, 42.35205, 41.7398, 40.78961, 
    39.63939, 38.49644, 37.53534, 56.86322, 56.48124, 56.29373,
  57.6715, 57.78593, 58.0331, 58.44473, 59.03896, 59.81201, 40.78123, 
    41.73415, 42.35238, 42.62211, 42.59517, 42.26209, 41.56049, 40.49372, 
    39.21342, 37.95061, 36.89904, 56.24854, 55.85274, 55.66045,
  56.71901, 56.85788, 57.15284, 57.63263, 58.31116, 59.181, 40.23441, 
    41.3254, 42.03205, 42.31787, 42.23014, 41.76385, 40.87186, 39.59026, 
    38.11946, 36.73368, 35.6408, 55.09318, 54.72622, 54.54812,
  55.57771, 55.73886, 56.07576, 56.61088, 57.35025, 58.27982, 39.36735, 
    40.5679, 41.35833, 41.6565, 41.48089, 40.82277, 39.66553, 38.11025, 
    36.43648, 34.96788, 33.91004, 53.51741, 53.21481, 53.06567,
  54.39848, 54.57779, 54.94736, 55.52066, 56.29176, 57.23478, 38.30464, 
    39.53991, 40.36725, 40.64995, 40.36061, 39.48266, 38.04605, 36.24118, 
    34.43232, 32.96629, 32.01558, 51.76559, 51.53625, 51.41926,
  53.31495, 53.50907, 53.90441, 54.50444, 55.28876, 56.21555, 37.24476, 
    38.42739, 39.21799, 39.43929, 39.02059, 37.94297, 36.29341, 34.34952, 
    32.52503, 31.14085, 30.315, 50.12937, 49.9495, 49.85439,
  52.40918, 52.61736, 53.03756, 53.664, 54.46165, 55.37103, 36.36428, 
    37.43113, 38.11755, 38.23591, 37.69394, 36.48318, 34.74205, 32.79772, 
    31.05487, 29.77566, 29.03224, 48.82079, 48.64961, 48.55883,
  51.70614, 51.93006, 52.37979, 53.04234, 53.86924, 54.78133, 35.75928, 
    36.68177, 37.22456, 37.21952, 36.58157, 35.32495, 33.61718, 31.78005, 
    30.16193, 28.96541, 28.24312, 47.91634, 47.71211, 47.60699,
  51.18284, 51.42145, 51.9011, 52.60786, 53.49006, 54.45216, 55.50565, 
    56.29232, 56.71482, 56.63289, 55.97269, 54.75881, 53.15021, 51.42387, 
    49.87104, 48.67282, 47.87974, 47.3047, 47.02905, 46.89749,
  50.84099, 51.09223, 51.5974, 52.34077, 53.26546, 54.26474, 55.32153, 
    56.0509, 56.41494, 56.29127, 55.61507, 54.41713, 52.85139, 51.17375, 
    49.65057, 48.45248, 47.6282, 46.95538, 46.62883, 46.4756,
  50.65107, 50.90972, 51.43042, 52.19754, 53.15225, 54.18245, 55.24451, 
    55.96439, 56.31336, 56.17565, 55.48811, 54.28176, 52.71121, 51.03243, 
    49.50898, 48.30698, 47.46949, 46.77003, 46.42208, 46.25954,
  54.1953, 54.40676, 54.82819, 55.43834, 56.18054, 56.9608, 57.64518, 
    58.16187, 58.36267, 58.18026, 57.59526, 56.64962, 55.45316, 54.16415, 
    52.94326, 51.90548, 51.1, 50.56414, 50.22325, 50.0667,
  54.47023, 54.6719, 55.07385, 55.65563, 56.36323, 57.10732, 57.76368, 
    58.26263, 58.46276, 58.29585, 57.7399, 56.83297, 55.67865, 54.42791, 
    53.23714, 52.22227, 51.43689, 50.91479, 50.58538, 50.43404,
  54.96231, 55.14825, 55.51986, 56.05993, 56.72018, 57.41843, 58.0439, 
    58.52871, 58.74001, 58.60577, 58.09747, 57.24561, 56.14559, 54.94141, 
    53.78746, 52.8036, 52.05031, 51.55366, 51.24416, 51.10123,
  55.63585, 55.80286, 56.13842, 56.63007, 57.23738, 57.88682, 58.47754, 
    58.95513, 59.18895, 59.10286, 58.66019, 57.88032, 56.84615, 55.69235, 
    54.5727, 53.6148, 52.88994, 52.42746, 52.13621, 51.99977,
  56.42105, 56.5699, 56.87083, 57.31653, 57.87466, 58.48119, 59.0281, 
    59.50849, 59.77232, 59.74407, 59.38207, 58.69164, 57.73548, 56.63225, 
    55.53443, 54.58182, 53.8618, 53.44377, 53.15785, 53.02113,
  57.21513, 57.35058, 57.62555, 58.03666, 58.55813, 59.13644, 59.63842, 
    60.13691, 60.43458, 60.46735, 60.19699, 59.61315, 58.74794, 57.69294, 
    56.59618, 55.61442, 54.85872, 54.47748, 54.17969, 54.03484,
  57.90846, 58.03843, 58.30169, 58.69539, 59.19502, 59.75664, 40.26481, 
    40.81186, 41.1501, 41.24372, 41.0743, 40.61882, 39.86699, 38.86784, 
    37.75817, 36.71462, 35.88257, 55.43645, 55.11127, 54.94825,
  58.37327, 58.5068, 58.77649, 59.17971, 59.69162, 60.2714, 40.89447, 
    41.45835, 41.806, 41.93946, 41.86703, 41.55555, 40.94879, 40.03872, 
    38.92756, 37.79944, 36.8419, 56.16454, 55.78291, 55.59231,
  58.53124, 58.67626, 58.96802, 59.40255, 59.95095, 60.56886, 41.28106, 
    41.85854, 42.20352, 42.34927, 42.32974, 42.11079, 41.60705, 40.7685, 
    39.66421, 38.4736, 37.4128, 56.57072, 56.13159, 55.91356,
  58.32774, 58.48969, 58.81497, 59.29838, 59.90658, 60.59002, 41.38776, 
    42.01425, 42.3767, 42.52566, 42.51624, 42.32112, 41.8439, 41.01426, 
    39.88333, 38.62699, 37.47732, 56.55905, 56.07699, 55.83973,
  57.74759, 57.9297, 58.29593, 58.84103, 59.52902, 60.30647, 41.2041, 
    41.93657, 42.35661, 42.51635, 42.48447, 42.24398, 41.70201, 40.78983, 
    39.564, 38.21214, 36.97928, 56.0644, 55.56473, 55.32148,
  56.82522, 57.02869, 57.43854, 58.04999, 58.82586, 59.71039, 40.71297, 
    41.5957, 42.11058, 42.2943, 42.21653, 41.86792, 41.16922, 40.0741, 
    38.67321, 37.19156, 35.89285, 55.06047, 54.5789, 54.34673,
  55.65211, 55.8759, 56.32637, 56.99754, 57.85013, 58.82547, 39.90641, 
    40.94014, 41.56249, 41.77624, 41.63424, 41.12672, 40.19454, 38.83466, 
    37.20314, 35.58784, 34.27322, 53.5969, 53.17244, 52.96843,
  54.36657, 54.60782, 55.09136, 55.80653, 56.70844, 57.7323, 38.83781, 
    39.96837, 40.67228, 40.90409, 40.68138, 39.9846, 38.78056, 37.1304, 
    35.27957, 33.58332, 32.32899, 51.84065, 51.49731, 51.33073,
  53.11951, 53.37517, 53.88384, 54.62668, 55.54894, 56.57557, 37.65399, 
    38.7911, 39.51442, 39.73075, 39.41375, 38.53082, 37.08196, 35.20462, 
    33.22921, 31.54478, 30.40713, 50.06146, 49.79034, 49.65609,
  52.03055, 52.29931, 52.82953, 53.59215, 54.51978, 55.52382, 36.54631, 
    37.60353, 38.27173, 38.42857, 38.01316, 36.98757, 35.38992, 33.42212, 
    31.45545, 29.85763, 28.83211, 48.52985, 48.29145, 48.17163,
  51.16138, 51.44458, 51.99934, 52.78629, 53.72396, 54.70736, 35.67949, 
    36.60775, 37.166, 37.22876, 36.72421, 35.6256, 34.00591, 32.0948, 
    30.24263, 28.7558, 27.79351, 47.41073, 47.1521, 47.02292,
  50.50953, 50.80715, 51.38917, 52.21203, 53.18808, 54.19568, 55.22095, 
    56.00345, 56.44391, 56.43165, 55.89485, 54.81758, 53.28255, 51.49911, 
    49.76013, 48.32147, 47.31913, 46.66538, 46.32566, 46.16497,
  50.0817, 50.39212, 50.99809, 51.85135, 52.85728, 53.88546, 54.92467, 
    55.64634, 56.03054, 55.9789, 55.42406, 54.35713, 52.8637, 51.14074, 
    49.45411, 48.037, 47.01506, 46.23205, 45.83475, 45.64887,
  49.84513, 50.16414, 50.78702, 51.66375, 52.69602, 53.74824, 54.79432, 
    55.50088, 55.86813, 55.8042, 55.24245, 54.17305, 52.68056, 50.96111, 
    49.27819, 47.86064, 46.82753, 46.00374, 45.58197, 45.38536,
  53.55328, 53.83249, 54.36798, 55.10173, 55.93909, 56.76576, 57.46073, 
    57.98362, 58.2277, 58.14237, 57.69647, 56.89129, 55.78012, 54.47587, 
    53.13298, 51.9043, 50.8978, 50.19124, 49.73436, 49.51944,
  53.89677, 54.16475, 54.67902, 55.38464, 56.19198, 56.99204, 57.66927, 
    58.18475, 58.43181, 58.35794, 57.93131, 57.15351, 56.07645, 54.80778, 
    53.49483, 52.2864, 51.29224, 50.59228, 50.13765, 49.92244,
  54.49146, 54.74477, 55.23209, 55.90353, 56.67614, 57.44664, 58.10382, 
    58.61479, 58.87166, 58.82032, 58.4275, 57.69294, 56.66372, 55.43898, 
    54.15815, 52.96811, 51.98442, 51.29439, 50.84108, 50.62418,
  55.26639, 55.50506, 55.96541, 56.60254, 57.33993, 58.07987, 58.70754, 
    59.21283, 59.4787, 59.4534, 59.10468, 58.42924, 57.46442, 56.2945, 
    55.047, 53.86741, 52.88126, 52.20321, 51.74271, 51.5194,
  56.12065, 56.34829, 56.7874, 57.39599, 58.10163, 58.81197, 59.39201, 
    59.88715, 60.15361, 60.1497, 59.84988, 59.24776, 58.36491, 57.26197, 
    56.04783, 54.86548, 53.85478, 53.1932, 52.71422, 52.47942,
  56.94144, 57.16372, 57.59064, 58.17957, 58.85911, 59.54282, 60.06839, 
    60.551, 60.80843, 60.81857, 60.5696, 60.05228, 59.26646, 58.23991, 
    57.0552, 55.851, 54.78798, 54.13115, 53.63059, 53.38403,
  57.63624, 57.85918, 58.28289, 58.85916, 59.51273, 60.16441, 40.70007, 
    41.18171, 41.42714, 41.44541, 41.25015, 40.83256, 40.16419, 39.22897, 
    38.07368, 36.82888, 35.68701, 54.94282, 54.43562, 54.18133,
  58.10994, 58.33978, 58.77208, 59.35169, 59.99759, 60.63238, 41.24575, 
    41.68703, 41.89892, 41.9199, 41.78304, 41.47444, 40.9369, 40.11306, 
    39.01091, 37.74379, 36.52636, 55.56274, 55.02207, 54.75021,
  58.31213, 58.55312, 59.00225, 59.59624, 60.24647, 60.87452, 41.53236, 
    41.94393, 42.13102, 42.15205, 42.05397, 41.81981, 41.37372, 40.63275, 
    39.57891, 38.30823, 37.043, 55.92801, 55.35035, 55.05944,
  58.20216, 58.45697, 58.92969, 59.5505, 60.22415, 60.87057, 41.56667, 
    41.98957, 42.18101, 42.20834, 42.12852, 41.92586, 41.51683, 40.80699, 
    39.76542, 38.47683, 37.16399, 55.97122, 55.36036, 55.05365,
  57.75655, 58.02706, 58.52982, 59.19194, 59.91364, 60.61243, 41.36634, 
    41.85596, 42.09002, 42.13605, 42.05783, 41.84432, 41.41314, 40.66946, 
    39.58158, 38.23442, 36.85421, 55.63802, 55.00314, 54.68705,
  56.97704, 57.26439, 57.80222, 58.51818, 59.30996, 60.09123, 40.92492, 
    41.52929, 41.83998, 41.91773, 41.82817, 41.56464, 41.05118, 40.20111, 
    38.99504, 37.53653, 36.06877, 54.88437, 54.24479, 53.93053,
  55.90461, 56.20857, 56.7825, 57.5564, 58.42665, 59.30161, 40.21576, 
    40.95647, 41.36303, 41.4811, 41.36976, 41.02203, 40.36933, 39.34006, 
    37.94381, 36.32933, 34.77707, 53.69593, 53.08371, 52.78742,
  54.62961, 54.94805, 55.55318, 56.37656, 57.31311, 58.26498, 39.22763, 
    40.08752, 40.58667, 40.74448, 40.60133, 40.14203, 39.30377, 38.03779, 
    36.40398, 34.62465, 33.03204, 52.12929, 51.58107, 51.31887,
  53.28505, 53.61446, 54.24149, 55.09616, 56.07051, 57.05979, 38.01597, 
    38.93836, 39.49879, 39.68056, 39.49343, 38.90692, 37.86441, 36.35087, 
    34.49493, 32.60248, 31.04608, 50.35303, 49.88869, 49.66716,
  52.01611, 52.35357, 52.99389, 53.86173, 54.84388, 55.82788, 36.72202, 
    37.62897, 38.19511, 38.36776, 38.12223, 37.41294, 36.19625, 34.50127, 
    32.52364, 30.6217, 29.16605, 48.63203, 48.23471, 48.04359,
  50.93852, 51.28405, 51.93573, 52.80959, 53.78395, 54.73743, 35.55392, 
    36.38323, 36.89742, 37.02043, 36.70366, 35.89832, 34.58519, 32.83835, 
    30.88861, 29.08304, 27.74526, 47.23436, 46.8499, 46.66276,
  50.10142, 50.45667, 51.12464, 52.01576, 53.00246, 53.95121, 54.80829, 
    55.5096, 55.93007, 55.9912, 55.63076, 54.80462, 53.51591, 51.85751, 
    50.04115, 48.35385, 47.05421, 46.27667, 45.81059, 45.58904,
  49.54, 49.90474, 50.58791, 51.49352, 52.48858, 53.43708, 54.34329, 
    54.99323, 55.36925, 55.39682, 55.01229, 54.17761, 52.90726, 51.29963, 
    49.55214, 47.92033, 46.63262, 45.68652, 45.16164, 44.91283,
  49.23097, 49.6046, 50.30347, 51.22738, 52.23906, 53.20028, 54.12563, 
    54.75952, 55.12002, 55.13682, 54.74604, 53.90971, 52.6427, 51.04288, 
    49.30492, 47.67902, 46.38522, 45.37478, 44.82244, 44.56149,
  53.56129, 53.85859, 54.41606, 55.15584, 55.9707, 56.74991, 57.3925, 
    57.88347, 58.137, 58.11073, 57.76998, 57.09885, 56.11912, 54.90449, 
    53.57964, 52.29543, 51.1881, 50.37351, 49.83055, 49.56888,
  53.91443, 54.2016, 54.74068, 55.45764, 56.25008, 57.01101, 57.64092, 
    58.12696, 58.38124, 58.36082, 58.03173, 57.37978, 56.42707, 55.24367, 
    53.94711, 52.68174, 51.5827, 50.7705, 50.22346, 49.95768,
  54.51342, 54.79013, 55.31057, 56.00497, 56.77558, 57.51827, 58.13164, 
    58.61262, 58.86885, 58.85885, 58.55058, 57.9308, 57.01876, 55.87616, 
    54.60998, 53.3582, 52.25865, 51.44673, 50.88882, 50.61462,
  55.27288, 55.54115, 56.04609, 56.72081, 57.47073, 58.19417, 58.77911, 
    59.25005, 59.50183, 59.49901, 59.21483, 58.63747, 57.7801, 56.69037, 
    55.45937, 54.21648, 53.10422, 52.29336, 51.71558, 51.42827,
  56.08652, 56.35006, 56.84481, 57.50402, 58.23403, 58.9362, 59.47499, 
    59.92888, 60.16549, 60.16134, 59.89965, 59.37115, 58.58022, 57.55488, 
    56.36425, 55.12539, 53.98668, 53.18136, 52.57851, 52.27631,
  56.85057, 57.11302, 57.6025, 58.24937, 58.95936, 59.63862, 60.12795, 
    60.56156, 60.77552, 60.76316, 60.52194, 60.04612, 59.32906, 58.37478, 
    57.22494, 55.98058, 54.79909, 53.98908, 53.36836, 53.05655,
  57.49243, 57.75611, 58.24226, 58.87474, 59.55672, 60.20265, 40.71272, 
    41.13792, 41.3306, 41.30607, 41.08488, 40.66875, 40.03691, 39.16242, 
    38.05218, 36.78643, 35.5413, 54.65519, 54.04969, 53.74195,
  57.93824, 58.20647, 58.69546, 59.32183, 59.98539, 60.60515, 41.18829, 
    41.57235, 41.73175, 41.69902, 41.50906, 41.1635, 40.62604, 39.84396, 
    38.79453, 37.53599, 36.2517, 55.17342, 54.55558, 54.24017,
  58.1512, 58.42612, 58.92199, 59.5475, 60.1981, 60.79621, 41.41687, 
    41.77092, 41.90857, 41.87365, 41.71065, 41.41962, 40.95225, 40.23977, 
    39.24214, 38.0016, 36.70021, 55.49062, 54.85296, 54.52605,
  58.09723, 58.38095, 58.88914, 59.52362, 60.17564, 60.76981, 41.41083, 
    41.76437, 41.90348, 41.87738, 41.73665, 41.48014, 41.05192, 40.37455, 
    39.39944, 38.15929, 36.83199, 55.55058, 54.88839, 54.54897,
  57.75069, 58.04588, 58.57397, 59.23212, 59.90742, 60.52423, 41.19263, 
    41.58464, 41.75369, 41.7501, 41.62788, 41.38529, 40.96285, 40.27949, 
    39.28375, 38.0057, 36.62289, 55.3054, 54.61616, 54.265,
  57.10047, 57.40968, 57.96553, 58.66305, 59.38507, 60.0524, 40.76386, 
    41.23093, 41.45589, 41.48692, 41.37837, 41.12775, 40.67487, 39.93847, 
    38.86899, 37.50364, 36.03096, 54.71071, 54, 53.64226,
  56.16189, 56.48627, 57.07439, 57.82143, 58.60616, 59.343, 40.10389, 
    40.66906, 40.96738, 41.04053, 40.93864, 40.65644, 40.13396, 39.29201, 
    38.08972, 36.58767, 35.0048, 53.73449, 53.02232, 52.66985,
  54.98978, 55.32782, 55.94614, 56.74134, 57.58897, 58.39569, 39.18939, 
    39.85273, 40.22878, 40.34507, 40.2401, 39.90168, 39.26898, 38.26785, 
    36.87786, 35.20686, 33.52778, 52.38423, 51.7045, 51.37403,
  53.68461, 54.03228, 54.67204, 55.5016, 56.39435, 57.2493, 38.03446, 
    38.76691, 39.20664, 39.35697, 39.23531, 38.8173, 38.04084, 36.84347, 
    35.24209, 33.41433, 31.69864, 50.75215, 50.13808, 49.84316,
  52.3807, 52.73341, 53.38345, 54.22768, 55.13763, 56.00527, 36.72802, 
    37.47573, 37.94363, 38.10439, 37.94739, 37.43391, 36.50508, 35.12255, 
    33.35465, 31.448, 29.78312, 49.04397, 48.50272, 48.24277,
  51.21339, 51.56926, 52.2233, 53.06837, 53.97211, 54.82025, 35.45986, 
    36.16963, 36.61963, 36.75528, 36.54111, 35.93038, 34.87872, 33.38579, 
    31.56999, 29.70831, 28.1675, 47.5403, 47.03501, 46.78886,
  50.27034, 50.63131, 51.29352, 52.14641, 53.05387, 53.89252, 54.57723, 
    55.18853, 55.57075, 55.65916, 55.39891, 54.74215, 53.66558, 52.20173, 
    50.48335, 48.7547, 47.31098, 46.45822, 45.88455, 45.60666,
  49.62043, 49.98686, 50.65652, 51.51394, 52.42045, 53.2534, 54.01965, 
    54.59556, 54.94751, 55.00941, 54.72148, 54.03977, 52.9542, 51.51268, 
    49.84961, 48.18636, 46.78065, 45.74793, 45.1265, 44.82475,
  49.26197, 49.6364, 50.31907, 51.18989, 52.10703, 52.94773, 53.7484, 
    54.31316, 54.65431, 54.70748, 54.41149, 53.7231, 52.63475, 51.19651, 
    49.54176, 47.88668, 46.47958, 45.36778, 44.72035, 44.40699,
  53.91416, 54.20295, 54.73398, 55.4199, 56.15446, 56.84116, 57.40083, 
    57.84185, 58.0922, 58.11541, 57.87584, 57.34785, 56.53111, 55.46394, 
    54.23191, 52.96254, 51.80058, 50.89743, 50.26821, 49.95542,
  54.24361, 54.52488, 55.04283, 55.7135, 56.43395, 57.10913, 57.65794, 
    58.09251, 58.33801, 58.35907, 58.1221, 57.60402, 56.80583, 55.76389, 
    54.55782, 53.30766, 52.15398, 51.25316, 50.61699, 50.29811,
  54.79301, 55.06955, 55.57914, 56.23975, 56.94988, 57.61469, 58.14651, 
    58.57106, 58.80733, 58.82411, 58.59221, 58.09177, 57.32316, 56.31607, 
    55.13932, 53.9033, 52.74652, 51.84306, 51.18966, 50.85862,
  55.47538, 55.75005, 56.2555, 56.90957, 57.61055, 58.2639, 58.76741, 
    59.17654, 59.39573, 59.4016, 59.17241, 58.69284, 57.96147, 56.99792, 
    55.85585, 54.63272, 53.46474, 52.56058, 51.88378, 51.53747,
  56.19242, 56.46725, 56.97083, 57.61892, 58.30885, 58.94809, 59.41126, 
    59.80088, 59.99576, 59.98325, 59.75197, 59.29268, 58.60187, 57.68724, 
    56.58415, 55.37371, 54.1889, 53.2892, 52.59129, 52.23187,
  56.85727, 57.13246, 57.63332, 58.27264, 58.94777, 59.57055, 59.99681, 
    60.36782, 60.53713, 60.50319, 60.26687, 59.8261, 59.17551, 58.31022, 
    57.24508, 56.042, 54.83194, 53.92823, 53.22363, 52.86062,
  57.41762, 57.6912, 58.18414, 58.80533, 59.45329, 60.04861, 40.5089, 
    40.87759, 41.02926, 40.97328, 40.72967, 40.30806, 39.70044, 38.88501, 
    37.85077, 36.63619, 35.37978, 54.42514, 53.7598, 53.41525,
  57.81677, 58.08929, 58.57565, 59.18121, 59.80566, 60.37596, 40.91454, 
    41.25608, 41.3851, 41.31685, 41.08161, 40.69305, 40.13821, 39.38294, 
    38.39798, 37.20295, 35.93579, 54.82481, 54.17031, 53.83006,
  58.02724, 58.29917, 58.77981, 59.37062, 59.97174, 60.51627, 41.09676, 
    41.41822, 41.53338, 41.46217, 41.24225, 40.88786, 40.37947, 39.6738, 
    38.73153, 37.56126, 36.29762, 55.0794, 54.4242, 54.08178,
  58.01957, 58.29296, 58.77243, 59.35536, 59.94152, 60.46867, 41.06134, 
    41.37712, 41.49232, 41.43058, 41.23405, 40.91464, 40.44497, 39.77404, 
    38.85676, 37.69558, 36.42117, 55.14075, 54.47167, 54.12144,
  57.76775, 58.04646, 58.5332, 59.12119, 59.70797, 60.23309, 40.82857, 
    41.15872, 41.29136, 41.25303, 41.08755, 40.80231, 40.36173, 39.70749, 
    38.78973, 37.60735, 36.28924, 54.96614, 54.26937, 53.90592,
  57.25357, 57.54212, 58.04631, 58.65523, 59.26212, 59.80465, 40.40584, 
    40.77205, 40.93933, 40.93594, 40.80461, 40.54723, 40.12097, 39.46035, 
    38.51015, 37.26804, 35.86703, 54.51455, 53.78166, 53.40281,
  56.4752, 56.77686, 57.30648, 57.94984, 58.59448, 59.17294, 39.78334, 
    40.20406, 40.41972, 40.45768, 40.3569, 40.11357, 39.67917, 38.98147, 
    37.96011, 36.61703, 35.10107, 53.74905, 52.98472, 52.59544,
  55.45797, 55.77291, 56.32996, 57.01308, 57.70446, 58.32951, 38.94112, 
    39.42534, 39.69686, 39.77693, 39.6967, 39.44594, 38.97167, 38.19649, 
    37.05924, 35.57899, 33.93961, 52.64985, 51.877, 51.49058,
  54.26565, 54.5905, 55.16934, 55.88627, 56.61986, 57.28785, 37.87367, 
    38.41365, 38.73822, 38.85435, 38.77909, 38.49338, 37.94083, 37.04374, 
    35.75154, 34.12081, 32.39132, 51.24883, 50.50319, 50.13649,
  53.00446, 53.33381, 53.92375, 54.65954, 55.41804, 56.10968, 36.62628, 
    37.19442, 37.55432, 37.6904, 37.59865, 37.24876, 36.584, 35.53703, 
    34.08604, 32.34254, 30.60488, 49.67531, 48.9848, 48.64729,
  51.80824, 52.13828, 52.73032, 53.46956, 54.23106, 54.91944, 35.34947, 
    35.91188, 36.27799, 36.40681, 36.27203, 35.83413, 35.04372, 33.86015, 
    32.30794, 30.55068, 28.91235, 48.17096, 47.52789, 47.20946,
  50.79364, 51.12561, 51.72179, 52.4669, 53.23347, 53.91843, 54.40244, 
    54.90225, 55.22894, 55.32751, 55.14959, 54.64972, 53.79424, 52.5777, 
    51.06141, 49.415, 47.91452, 47.01409, 46.3241, 45.9793,
  50.06843, 50.40219, 51.00018, 51.74516, 52.50947, 53.19145, 53.78865, 
    54.2743, 54.58864, 54.67056, 54.46391, 53.92426, 53.03004, 51.79608, 
    50.30027, 48.7079, 47.26465, 46.19009, 45.47517, 45.11524,
  49.66572, 50.00599, 50.61399, 51.36864, 52.14064, 52.82917, 53.4792, 
    53.96218, 54.27329, 54.35024, 54.13395, 53.58036, 52.6719, 51.42888, 
    49.9322, 48.34478, 46.90398, 45.73912, 45.0042, 44.63519,
  54.57228, 54.82514, 55.28344, 55.86408, 56.4743, 57.03749, 57.49353, 
    57.87067, 58.10467, 58.16346, 58.01218, 57.62106, 56.97657, 56.09066, 
    55.01101, 53.82915, 52.67648, 51.72601, 51.0268, 50.66648,
  54.8463, 55.09489, 55.54605, 56.1187, 56.72134, 57.27718, 57.72199, 
    58.0894, 58.31206, 58.3601, 58.20151, 57.80961, 57.17319, 56.30401, 
    55.24619, 54.08478, 52.94492, 52.00283, 51.30006, 50.93532,
  55.29827, 55.54727, 55.99865, 56.57055, 57.17023, 57.71976, 58.14568, 
    58.49754, 58.70055, 58.73021, 58.56014, 58.1685, 57.54591, 56.7007, 
    55.66867, 54.52474, 53.38778, 52.44949, 51.7328, 51.35754,
  55.85355, 56.1053, 56.56013, 57.13366, 57.73108, 58.27401, 58.67315, 
    59.00638, 59.18367, 59.18806, 59.00106, 58.60728, 57.99942, 57.18106, 
    56.17726, 55.05024, 53.91152, 52.9801, 52.2476, 51.86105,
  56.4323, 56.68634, 57.1431, 57.71558, 58.3079, 58.84338, 59.21193, 
    59.52768, 59.67776, 59.65311, 59.44455, 59.04442, 58.44826, 57.65523, 
    56.67915, 55.56807, 54.42544, 53.50442, 52.7639, 52.37135,
  56.96793, 57.22124, 57.6744, 58.23949, 58.82236, 59.3499, 59.69769, 
    60.00156, 60.12936, 60.07726, 59.84565, 59.43542, 58.84605, 58.0734, 
    57.12024, 56.01936, 54.86715, 53.94803, 53.21596, 52.82857,
  57.42582, 57.67304, 58.11245, 58.65695, 59.21715, 59.72741, 40.12022, 
    40.43256, 40.55144, 40.47447, 40.21726, 39.79391, 39.20802, 38.44929, 
    37.50521, 36.3899, 35.20277, 54.26243, 53.59024, 53.23577,
  57.76233, 58.00209, 58.42602, 58.94893, 59.48635, 59.97858, 40.45712, 
    40.75971, 40.86872, 40.77944, 40.5145, 40.094, 39.52331, 38.78939, 
    37.87167, 36.77254, 35.59061, 54.53179, 53.89172, 53.5539,
  57.95609, 58.18761, 58.59451, 59.0932, 59.60361, 60.07244, 40.60131, 
    40.89592, 40.99923, 40.90686, 40.64755, 40.24358, 39.69748, 38.99178, 
    38.10112, 37.02237, 35.85372, 54.7114, 54.08924, 53.75942,
  57.98111, 58.20607, 58.59891, 59.07648, 59.56177, 60.0068, 40.54622, 
    40.83394, 40.93657, 40.8526, 40.61488, 40.2434, 39.73312, 39.05914, 
    38.19154, 37.12395, 35.9534, 54.75989, 54.1356, 53.80391,
  57.81213, 58.03476, 58.42112, 58.88657, 59.35463, 59.78028, 40.30639, 
    40.59116, 40.70081, 40.63828, 40.43765, 40.11266, 39.64739, 39.00665, 
    38.15374, 37.07822, 35.87524, 54.63858, 53.98919, 53.64443,
  57.42785, 57.65379, 58.04415, 58.51058, 58.97412, 59.38986, 39.89206, 
    40.18149, 40.30744, 40.27719, 40.12319, 39.85094, 39.43296, 38.82206, 
    37.97128, 36.86327, 35.59147, 54.31076, 53.6159, 53.24861,
  56.81648, 57.05088, 57.4553, 57.93633, 58.41017, 58.82924, 39.30347, 
    39.60833, 39.75971, 39.76756, 39.66039, 39.43585, 39.05676, 38.46379, 
    37.59667, 36.42919, 35.05562, 53.74139, 52.99086, 52.59781,
  55.98264, 56.22812, 56.65263, 57.15802, 57.65483, 58.09085, 38.53048, 
    38.86156, 39.04581, 39.09204, 39.02264, 38.82859, 38.46619, 37.86589, 
    36.95457, 35.7003, 34.20676, 52.90027, 52.10164, 51.68926,
  54.9581, 55.21363, 55.65792, 56.19002, 56.71576, 57.17701, 37.56429, 
    37.92649, 38.14667, 38.22645, 38.17827, 37.98659, 37.60413, 36.95604, 
    35.96373, 34.60221, 33.00131, 51.78178, 50.96265, 50.54612,
  53.81401, 54.07558, 54.53341, 55.08633, 55.63705, 56.121, 36.42412, 
    36.81117, 37.06236, 37.16463, 37.11496, 36.88972, 36.44105, 35.69791, 
    34.59275, 33.12957, 31.48174, 50.4463, 49.64398, 49.23944,
  52.66398, 52.92748, 53.39103, 53.95419, 54.51722, 55.00991, 35.21988, 
    35.62035, 35.89048, 35.99675, 35.91771, 35.6214, 35.06378, 34.19118, 
    32.9706, 31.45679, 29.869, 49.06422, 48.30092, 47.91174,
  51.63531, 51.90114, 52.37117, 52.94558, 53.52117, 54.02063, 54.29196, 
    54.66435, 54.92081, 55.01367, 54.89964, 54.53778, 53.89389, 52.94442, 
    51.7003, 50.25198, 48.81049, 47.91793, 47.12893, 46.71832,
  50.86829, 51.13459, 51.60582, 52.18259, 52.76197, 53.26652, 53.6731, 
    54.0532, 54.3159, 54.40373, 54.26373, 53.85328, 53.14712, 52.14169, 
    50.87299, 49.44691, 48.06491, 47.01902, 46.23492, 45.8218,
  50.43756, 50.70901, 51.18842, 51.77404, 52.3621, 52.87532, 53.35176, 
    53.73924, 54.00779, 54.09599, 53.94638, 53.51569, 52.78262, 51.75121, 
    50.46501, 49.03319, 47.65383, 46.5119, 45.7179, 45.30001,
  55.9782, 56.13395, 56.41501, 56.76888, 57.13903, 57.48151, 57.75652, 
    58.01578, 58.1988, 58.27805, 58.22149, 57.99958, 57.5923, 56.99123, 
    56.2047, 55.27076, 54.27455, 53.38313, 52.66513, 52.27362,
  56.12603, 56.28106, 56.56086, 56.913, 57.28055, 57.61885, 57.88277, 
    58.13012, 58.29631, 58.35596, 58.27974, 58.0415, 57.62467, 57.02335, 
    56.24669, 55.33076, 54.35566, 53.4884, 52.78317, 52.39746,
  56.36995, 56.52831, 56.81278, 57.16852, 57.53653, 57.87128, 58.11709, 
    58.34643, 58.48553, 58.51333, 58.40586, 58.14287, 57.71265, 57.11116, 
    56.34574, 55.44711, 54.4882, 53.64454, 52.94656, 52.56329,
  56.67311, 56.8353, 57.12505, 57.48494, 57.85432, 58.18761, 58.41399, 
    58.62637, 58.7361, 58.72702, 58.58193, 58.28802, 57.83926, 57.23354, 
    56.47578, 55.5904, 54.64304, 53.82343, 53.13461, 52.75536,
  56.99488, 57.15829, 57.44926, 57.80983, 58.17984, 58.51476, 58.72806, 
    58.92981, 59.01488, 58.9705, 58.78655, 58.45817, 57.98548, 57.36896, 
    56.61193, 55.73317, 54.79217, 53.99123, 53.31927, 52.94966,
  57.30004, 57.46011, 57.74545, 58.10099, 58.47005, 58.80936, 59.02379, 
    59.22347, 59.29349, 59.22029, 58.99998, 58.63552, 58.13364, 57.49864, 
    56.73358, 55.85247, 54.91067, 54.11666, 53.47119, 53.11897,
  57.57504, 57.7248, 57.99277, 58.33018, 58.68731, 59.02438, 39.2887, 
    39.50799, 39.58018, 39.48415, 39.22652, 38.82185, 38.28339, 37.61689, 
    36.82206, 35.90628, 34.93155, 54.15247, 53.57986, 53.27415,
  57.79063, 57.92786, 58.17518, 58.4911, 58.83265, 59.16311, 39.51643, 
    39.74436, 39.82071, 39.71542, 39.43834, 39.00922, 38.44628, 37.75977, 
    36.95194, 36.0303, 35.06362, 54.21628, 53.6947, 53.41879,
  57.93076, 58.05314, 58.27524, 58.56282, 58.87962, 59.19342, 39.6065, 
    39.83959, 39.91884, 39.81091, 39.53013, 39.09883, 38.535, 37.84835, 
    37.04145, 36.12304, 35.16886, 54.26715, 53.78365, 53.52834,
  57.97306, 58.08029, 58.2759, 58.53178, 58.81764, 59.10577, 39.53246, 
    39.76011, 39.83841, 39.73568, 39.4702, 39.06306, 38.52628, 37.86308, 
    37.0722, 36.16158, 35.21067, 54.27351, 53.80413, 53.55621,
  57.89428, 57.98846, 58.16032, 58.38564, 58.63835, 58.89423, 39.29821, 
    39.5097, 39.58503, 39.49729, 39.2665, 38.90844, 38.42453, 37.80647, 
    37.04408, 36.14004, 35.17271, 54.20122, 53.71691, 53.46019,
  57.67295, 57.75832, 57.9129, 58.1134, 58.33554, 58.55701, 38.91313, 
    39.10105, 39.17355, 39.10964, 38.92809, 38.6366, 38.22402, 37.6675, 
    36.94286, 36.0411, 35.03342, 54.01907, 53.4903, 53.20825,
  57.29232, 57.3742, 57.52024, 57.70514, 57.90392, 58.09457, 38.38602, 
    38.5489, 38.62067, 38.58561, 38.4588, 38.23945, 37.90495, 37.41756, 
    36.7351, 35.8302, 34.76004, 53.69926, 53.10162, 52.78109,
  56.74211, 56.82553, 56.97195, 57.15199, 57.33818, 57.50747, 37.72108, 
    37.86424, 37.93919, 37.93325, 37.85622, 37.7003, 37.43499, 37.01019, 
    36.36484, 35.44945, 34.30256, 53.214, 52.53499, 52.17054,
  56.02409, 56.11262, 56.2665, 56.45182, 56.63768, 56.7989, 36.91954, 
    37.05321, 37.1364, 37.156, 37.11462, 36.99909, 36.77537, 36.38642, 
    35.75717, 34.82013, 33.59835, 52.53863, 51.78457, 51.38153,
  55.16484, 55.25997, 55.42531, 55.62328, 55.81905, 55.98453, 35.99166, 
    36.12795, 36.22481, 36.26381, 36.23724, 36.12659, 35.89798, 35.49531, 
    34.84218, 33.87022, 32.60382, 51.67203, 50.87105, 50.44451,
  54.23248, 54.33412, 54.51184, 54.72521, 54.93483, 55.10965, 35.00769, 
    35.16297, 35.28099, 35.33203, 35.29546, 35.14672, 34.85426, 34.37194, 
    33.64181, 32.62506, 31.37923, 50.67691, 49.87352, 49.44065,
  53.33402, 53.44398, 53.63821, 53.87345, 54.10337, 54.29215, 54.25208, 
    54.41686, 54.54823, 54.60723, 54.55541, 54.35808, 53.98729, 53.41611, 
    52.62205, 51.61254, 50.47778, 49.75601, 48.94061, 48.48625,
  52.62133, 52.73528, 52.93833, 53.18711, 53.43276, 53.63625, 53.73211, 
    53.92769, 54.0866, 54.15733, 54.09124, 53.84931, 53.40726, 52.75166, 
    51.884, 50.84146, 49.73782, 48.9065, 48.12938, 47.68808,
  52.21372, 52.33232, 52.54416, 52.80486, 53.0638, 53.27942, 53.45597, 
    53.67013, 53.84631, 53.92611, 53.85511, 53.59183, 53.11391, 52.41455, 
    51.5055, 50.43502, 49.32563, 48.40167, 47.62848, 47.18734,
  57.05767, 57.13149, 57.26844, 57.44641, 57.63837, 57.82189, 57.96639, 
    58.13578, 58.26833, 58.33815, 58.31517, 58.17245, 57.8919, 57.46268, 
    56.88187, 56.16397, 55.36155, 54.61701, 53.9798, 53.6206,
  57.10897, 57.18298, 57.32003, 57.49773, 57.68869, 57.87014, 58.00613, 
    58.16563, 58.28219, 58.33125, 58.28485, 58.11922, 57.81987, 57.37949, 
    56.79804, 56.09133, 55.30994, 54.59618, 53.98316, 53.63812,
  57.19683, 57.27297, 57.41285, 57.59264, 57.78403, 57.96412, 58.08641, 
    58.23116, 58.32211, 58.33745, 58.25362, 58.05254, 57.72536, 57.2688, 
    56.68473, 55.98802, 55.22514, 54.54388, 53.95357, 53.62173,
  57.31436, 57.39238, 57.5348, 57.71695, 57.91026, 58.09202, 58.20218, 
    58.33408, 58.39814, 58.37542, 58.24799, 58.00481, 57.64338, 57.1646, 
    56.57199, 55.87905, 55.12846, 54.47614, 53.90985, 53.59253,
  57.44962, 57.52747, 57.66964, 57.85257, 58.04911, 58.23693, 58.34434, 
    58.46957, 58.51213, 58.4543, 58.28393, 57.9971, 57.59748, 57.09028, 
    56.48114, 55.78305, 55.03657, 54.40046, 53.86099, 53.56091,
  57.58821, 57.6627, 57.80022, 57.98105, 58.18143, 58.37886, 58.49714, 
    58.62285, 58.65316, 58.5677, 58.35892, 58.02935, 57.58844, 57.04621, 
    56.41166, 55.69882, 54.94844, 54.31441, 53.80342, 53.5233,
  57.72866, 57.79375, 57.9166, 58.08432, 58.27956, 58.48104, 38.64384, 
    38.7893, 38.82463, 38.71877, 38.47226, 38.09681, 37.60682, 37.01443, 
    36.32952, 35.56679, 34.77892, 54.17249, 53.72754, 53.49329,
  57.84931, 57.90309, 58.00817, 58.15894, 58.34395, 58.54316, 38.78834, 
    38.94623, 38.98957, 38.87644, 38.60851, 38.20078, 37.67178, 37.03937, 
    36.31982, 35.53449, 34.74888, 54.10058, 53.70694, 53.50406,
  57.93601, 57.97523, 58.05632, 58.18133, 58.34512, 58.53086, 38.83661, 
    39.0031, 39.05195, 38.93649, 38.66159, 38.24413, 37.70268, 37.0557, 
    36.32183, 35.52706, 34.74833, 54.06007, 53.70967, 53.53129,
  57.9676, 57.99013, 58.04282, 58.13514, 58.26836, 58.42946, 38.75139, 
    38.91359, 38.96147, 38.84885, 38.58411, 38.18353, 37.66114, 37.03018, 
    36.30611, 35.51521, 34.74063, 54.02598, 53.69769, 53.5315,
  57.92205, 57.92757, 57.95049, 58.00658, 58.10282, 58.22967, 38.52956, 
    38.67295, 38.7144, 38.61164, 38.37498, 38.01704, 37.54342, 36.95707, 
    36.2646, 35.48656, 34.70567, 53.96694, 53.63375, 53.46407,
  57.77957, 57.76989, 57.7653, 57.78592, 57.84293, 57.92929, 38.17734, 
    38.28921, 38.32041, 38.23424, 38.04036, 37.74514, 37.34358, 36.82529, 
    36.18282, 35.42402, 34.62309, 53.85438, 53.48774, 53.29763,
  57.52477, 57.5035, 57.47695, 57.46702, 57.48722, 57.53175, 37.70471, 
    37.7773, 37.79636, 37.73088, 37.58742, 37.36504, 37.04848, 36.61341, 
    36.0347, 35.30051, 34.46734, 53.66535, 53.23917, 53.01328,
  57.14633, 57.11818, 57.07745, 57.04538, 57.03589, 57.04343, 37.12193, 
    37.15511, 37.16273, 37.11839, 37.02384, 36.8715, 36.63849, 36.28876, 
    35.77885, 35.07274, 34.20081, 53.37859, 52.87412, 52.60207,
  56.63895, 56.60899, 56.56301, 56.51973, 56.49187, 56.47352, 36.43941, 
    36.44157, 36.44177, 36.41617, 36.36021, 36.26106, 36.09209, 35.81057, 
    35.35885, 34.67852, 33.77113, 52.97266, 52.38441, 52.06429,
  56.01256, 55.98546, 55.94305, 55.90039, 55.86742, 55.8377, 35.67379, 
    35.66175, 35.66283, 35.65271, 35.6185, 35.54263, 35.39846, 35.14361, 
    34.7166, 34.04935, 33.12514, 52.43378, 51.77622, 51.41667,
  55.30866, 55.28808, 55.25634, 55.22396, 55.1963, 55.16673, 34.88432, 
    34.88589, 34.90362, 34.9078, 34.87569, 34.78474, 34.61026, 34.31713, 
    33.85532, 33.17247, 32.26545, 51.77838, 51.09263, 50.71165,
  54.60598, 54.59632, 54.58385, 54.57324, 54.56156, 54.54022, 54.31188, 
    54.33621, 54.37673, 54.39944, 54.36792, 54.25018, 54.02285, 53.66381, 
    53.14848, 52.4612, 51.63381, 51.13912, 50.439, 50.03256,
  54.03268, 54.0298, 54.03039, 54.03685, 54.04163, 54.03239, 53.91666, 
    53.97623, 54.05069, 54.09364, 54.05936, 53.91102, 53.62634, 53.19155, 
    52.59951, 51.86144, 51.04162, 50.46848, 49.80909, 49.41685,
  53.70453, 53.70602, 53.71533, 53.73383, 53.75116, 53.7514, 53.70856, 
    53.78791, 53.88274, 53.9392, 53.90583, 53.74276, 53.42808, 52.95226, 
    52.31651, 51.54378, 50.71251, 50.0587, 49.4047, 49.01098 ;

 hu =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -0.1106728, -1.424353, -4.358764, -4.531942, -1.615602, 
    -0.1287433, 0, 0, 0, 0, 0, 0.1287433, 1.615602, 4.531942, 4.358764, 
    1.424353, 0.1106728,
  0, 0, 0, -1.988207, -11.85714, -28.03266, -28.77494, -12.98619, -2.243248, 
    0, 0, 0, 0, 0, 2.243248, 12.98619, 28.77494, 28.03266, 11.85714, 1.988207,
  0, 0, 0, -10.58723, -64.99364, -144.3692, -130.2805, -46.59549, -7.613373, 
    0, 0, 0, 0, 0, 7.613373, 46.59549, 130.2804, 144.3692, 64.99364, 10.58723,
  0, 0, 0, -12.64522, -77.50148, -171.5085, -154.8044, -58.58395, -10.18297, 
    0, 0, 0, 0, 0, 10.18297, 58.58395, 154.8044, 171.5085, 77.50148, 12.64522,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.76649, -79.25483, -176.0672, -159.1111, -60.7706, -10.58736, 
    0, 0, 0, 0, 0, 10.58736, 60.7706, 159.1111, 176.0672, 79.25483, 12.76649,
  0, 0, 0, -12.64522, -77.50148, -171.5085, -154.8044, -58.58395, -10.18297, 
    0, 0, 0, 0, 0, 10.18297, 58.58395, 154.8044, 171.5085, 77.50148, 12.64522,
  0, 0, 0, -10.58723, -64.99364, -144.3692, -130.2805, -46.59549, -7.613373, 
    0, 0, 0, 0, 0, 7.613373, 46.59549, 130.2804, 144.3692, 64.99364, 10.58723,
  0, 0, 0, -1.988207, -11.85714, -28.03266, -28.77494, -12.98619, -2.243248, 
    0, 0, 0, 0, 0, 2.243248, 12.98619, 28.77494, 28.03266, 11.85714, 1.988207,
  0, 0, 0, -0.1106728, -1.424353, -4.358764, -4.531942, -1.615602, 
    -0.1287433, 0, 0, 0, 0, 0, 0.1287433, 1.615602, 4.531942, 4.358764, 
    1.424353, 0.1106728,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -9.645885e-05, -0.003138623, -0.03697342, -0.1972138, -0.471016, 
    -0.4951233, -0.2278209, -0.04405944, -0.003739635, -0.0001112987, 0, 
    0.0001112987, 0.003739635, 0.04405944, 0.2278209, 0.4951233, 0.471016, 
    0.19711, 0.03382738,
  0, -0.003644529, -0.07429843, -0.5720896, -2.28144, -4.850519, -5.129148, 
    -2.667596, -0.6936634, -0.09125484, -0.004454046, 0, 0.004454046, 
    0.09125484, 0.6936634, 2.667596, 5.129148, 4.850519, 2.277797, 0.4977923,
  0, -0.05175889, -0.6866534, -3.80572, -11.51663, -20.77404, -21.66175, 
    -12.90584, -4.394247, -0.8121275, -0.06367584, 0, 0.06367584, 0.8121275, 
    4.394247, 12.90584, 21.66175, 20.77404, 11.46483, 3.119064,
  0, -0.3510744, -3.521681, -14.78139, -34.24212, -50.94402, -52.3101, 
    -36.21666, -15.63128, -3.765846, -0.3849536, 0, 0.3849536, 3.765846, 
    15.63128, 36.21666, 52.3101, 50.94402, 33.89231, 11.26234,
  0, -1.116555, -11.39667, -48.34528, -108.8036, -149.0275, -133.5865, 
    -75.27055, -29.9594, -6.956295, -0.6862993, 0, 0.6862993, 6.956295, 
    29.9594, 75.27055, 133.5865, 149.0274, 107.727, 37.00165,
  0, -1.433281, -14.64716, -61.83953, -137.0734, -187.2945, -168.4538, 
    -98.06427, -40.91406, -9.996977, -1.038464, 0, 1.038464, 9.996977, 
    40.91406, 98.06427, 168.4538, 187.2945, 135.7011, 47.27648,
  0, -1.485358, -15.38204, -65.96331, -148.0887, -203.6059, -183.1557, 
    -107.7188, -45.4556, -11.26227, -1.19079, 0, 1.19079, 11.26227, 45.4556, 
    107.7188, 183.1557, 203.6059, 146.6678, 50.67165,
  0, -1.489202, -15.46767, -66.66711, -150.6115, -207.284, -186.5588, 
    -110.1894, -46.61765, -11.57875, -1.228485, 0, 1.228485, 11.57875, 
    46.61765, 110.1894, 186.5588, 207.284, 149.187, 51.29039,
  0, -1.489306, -15.47138, -66.71632, -150.8723, -207.6383, -186.9032, 
    -110.474, -46.75299, -11.61462, -1.232733, 0, 1.232733, 11.61462, 
    46.75299, 110.474, 186.9032, 207.6383, 149.4477, 51.3359,
  0, -1.489306, -15.47138, -66.71632, -150.8723, -207.6383, -186.9032, 
    -110.474, -46.75299, -11.61462, -1.232733, 0, 1.232733, 11.61462, 
    46.75299, 110.474, 186.9032, 207.6383, 149.4477, 51.3359,
  0, -1.489306, -15.47138, -66.71632, -150.8723, -207.6383, -186.9032, 
    -110.474, -46.75299, -11.61462, -1.232733, 0, 1.232733, 11.61462, 
    46.75299, 110.474, 186.9032, 207.6383, 149.4477, 51.3359,
  0, -1.489202, -15.46767, -66.66711, -150.6115, -207.284, -186.5588, 
    -110.1894, -46.61765, -11.57875, -1.228485, 0, 1.228485, 11.57875, 
    46.61765, 110.1894, 186.5588, 207.284, 149.187, 51.29039,
  0, -1.485358, -15.38204, -65.96331, -148.0887, -203.6059, -183.1557, 
    -107.7188, -45.4556, -11.26227, -1.19079, 0, 1.19079, 11.26227, 45.4556, 
    107.7188, 183.1557, 203.6059, 146.6678, 50.67165,
  0, -1.433281, -14.64716, -61.83953, -137.0734, -187.2945, -168.4538, 
    -98.06427, -40.91406, -9.996977, -1.038464, 0, 1.038464, 9.996977, 
    40.91406, 98.06427, 168.4538, 187.2945, 135.7011, 47.27648,
  0, -1.116555, -11.39667, -48.34528, -108.8036, -149.0275, -133.5865, 
    -75.27055, -29.9594, -6.956295, -0.6862993, 0, 0.6862993, 6.956295, 
    29.9594, 75.27055, 133.5865, 149.0274, 107.727, 37.00165,
  0, -0.3510744, -3.521681, -14.78139, -34.24212, -50.94402, -52.3101, 
    -36.21666, -15.63126, -3.765846, -0.3849684, 0, 0.3849684, 3.765846, 
    15.63126, 36.21666, 52.3101, 50.94402, 33.89231, 11.26234,
  0, -0.05175889, -0.6866534, -3.80572, -11.51663, -20.77404, -21.66175, 
    -12.90584, -4.394247, -0.8121275, -0.06367584, 0, 0.06367584, 0.8121275, 
    4.394247, 12.90584, 21.66175, 20.77404, 11.46483, 3.119064,
  0, -0.003644529, -0.07544857, -0.5975122, -2.467687, -5.357205, -5.670953, 
    -2.897055, -0.727339, -0.09299534, -0.004470198, 0, 0.004470198, 
    0.09299534, 0.727339, 2.897055, 5.670953, 5.357205, 2.464058, 0.5220798,
  0, -7.915459e-05, -0.0009498551, -0.006181254, -0.02308436, -0.04674438, 
    -0.04880241, -0.02607065, -0.007275026, -0.001129752, -9.354635e-05, 0, 
    9.354635e-05, 0.001129752, 0.007275026, 0.02607065, 0.04880241, 
    0.04674438, 0.02299801, 0.005224204,
  -0.0001545453, -0.002564055, -0.02183284, -0.1114434, -0.3564464, 
    -0.6823246, -0.7216957, -0.4159781, -0.1363909, -0.02724493, 
    -0.003212442, 0, 0.003212442, 0.02724493, 0.1363909, 0.4159781, 
    0.7216957, 0.6821702, 0.353868, 0.08959621,
  -0.002769891, -0.03361034, -0.219796, -0.9036537, -2.467294, -4.387971, 
    -4.678451, -2.932265, -1.129686, -0.2813469, -0.0433618, 0, 0.0433618, 
    0.2813469, 1.129686, 2.932265, 4.678327, 4.385085, 2.433637, 0.6838038,
  -0.02634797, -0.2498512, -1.300066, -4.37655, -10.09203, -16.18374, 
    -17.14941, -11.74054, -5.308165, -1.616383, -0.3163989, 0, 0.3163989, 
    1.616383, 5.308165, 11.74054, 17.14806, 16.15567, 9.840928, 3.075615,
  -0.1552197, -1.203995, -5.136436, -14.24027, -27.21746, -37.98634, 
    -39.54972, -29.84263, -15.79911, -5.78855, -1.388415, 0, 1.388415, 
    5.78855, 15.79911, 29.84263, 39.5394, 37.81916, 26.00781, 9.099982,
  -0.6042287, -4.083549, -14.74194, -33.79564, -53.14474, -64.03078, 
    -66.48439, -56.11797, -34.39825, -14.71431, -4.084993, 0, 4.084993, 
    14.71431, 34.39825, 56.11797, 66.44025, 63.38972, 49.08347, 19.07141,
  -1.506048, -10.22478, -36.97513, -83.40836, -125.8726, -140.9819, 
    -128.2147, -89.97349, -50.08894, -20.38713, -5.453694, 0, 5.453694, 
    20.38713, 50.08894, 89.97349, 128.1389, 139.5529, 116.1764, 46.81511,
  -1.997113, -13.57499, -48.86349, -108.3481, -160.2497, -180.8471, 
    -166.4043, -118.6279, -68.03322, -28.71218, -7.991757, 0, 7.991757, 
    28.71218, 68.03322, 118.6279, 166.3092, 178.9995, 147.5378, 60.12846,
  -2.144811, -14.75771, -53.89066, -120.8711, -180.0647, -205.1317, 
    -188.7007, -134.848, -78.12237, -33.47867, -9.506922, 0, 9.506922, 
    33.47867, 78.12237, 134.848, 188.6, 203.1562, 166.2827, 67.72356,
  -2.172295, -15.03328, -55.35542, -125.329, -188.186, -214.7549, -197.5023, 
    -141.7438, -82.49405, -35.54688, -10.1664, 0, 10.1664, 35.54688, 
    82.49405, 141.7438, 197.3994, 212.7512, 174.1472, 70.73805,
  -2.17533, -15.07321, -55.6314, -126.392, -190.4884, -217.297, -199.8781, 
    -143.8313, -83.84976, -36.18324, -10.36676, 0, 10.36676, 36.18324, 
    83.84976, 143.8313, 199.7743, 215.2883, 176.4108, 71.52785,
  -2.175502, -15.07629, -55.65977, -126.5325, -190.8521, -217.6587, -200.227, 
    -144.1801, -84.08284, -36.29219, -10.40066, 0, 10.40066, 36.29219, 
    84.08284, 144.1801, 200.1231, 215.6494, 176.7713, 71.6403,
  -2.17533, -15.07321, -55.6314, -126.392, -190.4884, -217.297, -199.8781, 
    -143.8313, -83.84976, -36.18324, -10.36676, 0, 10.36676, 36.18324, 
    83.84976, 143.8313, 199.7743, 215.2883, 176.4108, 71.52785,
  -2.172295, -15.03328, -55.35542, -125.329, -188.186, -214.7549, -197.5023, 
    -141.7438, -82.49405, -35.54688, -10.1664, 0, 10.1664, 35.54688, 
    82.49405, 141.7438, 197.3994, 212.7512, 174.1472, 70.73805,
  -2.144811, -14.75771, -53.89066, -120.8711, -180.0647, -205.1317, 
    -188.7007, -134.848, -78.12237, -33.47867, -9.506922, 0, 9.506922, 
    33.47867, 78.12237, 134.848, 188.6, 203.1562, 166.2827, 67.72356,
  -1.997113, -13.57499, -48.86349, -108.3481, -160.2497, -180.8471, 
    -166.4043, -118.6279, -68.03322, -28.71218, -7.991757, 0, 7.991757, 
    28.71218, 68.03322, 118.6279, 166.3092, 178.9995, 147.5378, 60.12846,
  -1.506048, -10.22478, -36.97513, -83.40836, -125.8726, -140.9819, 
    -128.2147, -89.97348, -50.08894, -20.38713, -5.453707, 0, 5.453707, 
    20.38713, 50.08894, 89.97348, 128.1389, 139.5529, 116.1764, 46.81511,
  -0.6042287, -4.083579, -14.74259, -33.80119, -53.16919, -64.08242, 
    -66.53701, -56.14617, -34.40788, -14.71722, -4.085834, 0, 4.085834, 
    14.71722, 34.40788, 56.14617, 66.49287, 63.44136, 49.1079, 19.07632,
  -0.1552532, -1.205235, -5.151745, -14.33966, -27.59096, -38.76148, 
    -40.38325, -30.3223, -15.96086, -5.825705, -1.394756, 0, 1.394756, 
    5.825705, 15.96086, 30.3223, 40.37291, 38.59425, 26.38007, 9.184065,
  -0.02713067, -0.2672406, -1.458261, -5.176821, -12.60561, -21.03816, 
    -22.43792, -14.97079, -6.464798, -1.871175, -0.3489468, 0, 0.3489468, 
    1.871175, 6.464798, 14.97079, 22.43656, 21.00931, 12.33709, 3.717647,
  -0.007686974, -0.04793812, -0.1908363, -0.5645118, -1.244568, -1.973971, 
    -2.104207, -1.480072, -0.7163503, -0.2510944, -0.06300731, 0, 0.06300731, 
    0.2510944, 0.7163337, 1.479965, 2.103072, 1.965065, 1.196353, 0.3735716,
  -0.04870551, -0.2613763, -0.8819612, -2.250473, -4.416636, -6.585798, 
    -7.061854, -5.317093, -2.892844, -1.177021, -0.346752, 0, 0.346752, 
    1.177019, 2.89276, 5.316066, 7.052461, 6.52683, 4.152205, 1.367271,
  -0.2355841, -1.123383, -3.304671, -7.414326, -13.02617, -18.10315, 
    -19.30803, -15.37519, -9.22263, -4.243443, -1.423617, 0, 1.423617, 
    4.243422, 9.222062, 15.368, 19.25213, 17.80574, 11.88151, 4.100965,
  -0.8577683, -3.677983, -9.467377, -18.55865, -28.74956, -36.5085, 
    -38.42647, -32.41272, -21.3901, -11.0504, -4.166743, 0, 4.166743, 
    11.05025, 21.38688, 32.37738, 38.18594, 35.38828, 24.9827, 9.05652,
  -2.437775, -9.505665, -21.4459, -36.40242, -49.09857, -56.39412, -58.91578, 
    -53.21884, -38.63484, -22.18379, -9.230819, 0, 9.230819, 22.1832, 
    38.62237, 53.09417, 58.14224, 53.14919, 39.3769, 14.8865,
  -5.620964, -20.18425, -40.09894, -58.89241, -69.51617, -73.05064, 
    -77.29076, -75.80077, -60.35648, -37.90912, -17.00006, 0, 17.00006, 
    37.9077, 60.32531, 75.48383, 75.37769, 65.56701, 49.09581, 18.79547,
  -11.23946, -40.04322, -78.07516, -111.6943, -127.5791, -125.9439, 
    -117.1216, -98.12746, -70.63226, -41.87642, -18.17212, 0, 18.17212, 
    41.87554, 70.60988, 97.83334, 114.3433, 112.5407, 89.2264, 34.75319,
  -15.13974, -53.50325, -102.2562, -142.6409, -160.9448, -162.4527, 
    -154.7088, -130.3726, -94.77353, -57.01437, -25.16153, 0, 25.16153, 
    57.01338, 94.74815, 130.0298, 151.2063, 144.9267, 110.4985, 42.3222,
  -17.25249, -61.39297, -117.9381, -164.7632, -186.7229, -191.8679, 
    -183.1934, -152.9296, -111.3324, -67.54559, -30.15845, 0, 30.15845, 
    67.54446, 111.3045, 152.5632, 179.3672, 172.1876, 129.202, 49.25211,
  -18.12402, -64.99889, -126.0439, -177.4393, -202.2766, -208.9548, 
    -199.2558, -166.021, -121.182, -73.91232, -33.2123, 0, 33.2123, 73.91103, 
    121.1515, 165.6329, 195.2729, 188.3517, 141.446, 54.0176,
  -18.39265, -66.25471, -129.3021, -183.1927, -209.8062, -216.7003, 
    -206.4942, -172.3764, -126.1124, -77.12579, -34.75288, 0, 34.75288, 
    77.1244, 126.08, 171.9728, 202.4337, 195.7789, 147.7794, 56.56323,
  -18.44394, -66.5229, -130.0888, -184.728, -211.927, -218.7523, -208.4222, 
    -174.1963, -127.5582, -78.072, -35.2052, 0, 35.2052, 78.07059, 127.5251, 
    173.7871, 204.3376, 197.7606, 149.6358, 57.31929,
  -18.39265, -66.25471, -129.3021, -183.1927, -209.8062, -216.7003, 
    -206.4942, -172.3764, -126.1124, -77.12579, -34.75288, 0, 34.75288, 
    77.1244, 126.08, 171.9728, 202.4337, 195.7789, 147.7794, 56.56323,
  -18.12402, -64.99889, -126.0439, -177.4393, -202.2766, -208.9548, 
    -199.2558, -166.021, -121.182, -73.91232, -33.2123, 0, 33.2123, 73.91103, 
    121.1515, 165.6329, 195.2729, 188.3517, 141.446, 54.0176,
  -17.25249, -61.39297, -117.9382, -164.7636, -186.7237, -191.8683, 
    -183.1935, -152.9298, -111.3326, -67.54576, -30.15854, 0, 30.15854, 
    67.54463, 111.3047, 152.5635, 179.3673, 172.188, 129.2028, 49.25235,
  -15.13976, -53.50355, -102.2581, -142.6484, -160.9624, -162.4692, 
    -154.7187, -130.3797, -94.77895, -57.01835, -25.16368, 0, 25.16368, 
    57.01736, 94.75357, 130.0368, 151.2159, 144.9431, 110.516, 42.32787,
  -11.23997, -40.04755, -78.09814, -111.7748, -127.7636, -126.187, -117.3133, 
    -98.24487, -70.70638, -41.92001, -18.19234, 0, 18.19234, 41.91912, 
    70.68394, 97.95013, 114.5337, 112.7833, 89.40767, 34.81132,
  -5.625929, -20.22054, -40.26419, -59.41638, -70.68903, -74.88341, 
    -79.18588, -77.13098, -61.0724, -38.23548, -17.12114, 0, 17.12114, 
    38.23403, 61.04099, 76.81277, 77.27016, 67.39383, 50.2339, 19.15508,
  -2.47102, -9.715372, -22.27203, -38.75493, -54.01585, -63.92157, -67.02145, 
    -59.34806, -42.07701, -23.69606, -9.732143, 0, 9.732143, 23.69544, 
    42.06424, 59.22156, 66.24055, 60.63689, 44.0841, 16.41319,
  -1.018951, -4.566019, -12.4856, -26.12541, -43.08136, -57.32081, -61.04583, 
    -50.44147, -32.07829, -15.85297, -5.723922, 0, 5.723922, 15.85283, 
    32.07481, 50.40277, 60.77501, 56.00402, 38.41095, 13.59768,
  -0.2276659, -0.9316174, -2.367013, -4.849323, -8.167625, -11.21236, 
    -12.07136, -9.967039, -6.416276, -3.285159, -1.254022, -3.31091e-06, 
    1.253968, 3.284791, 6.413361, 9.94906, 11.98629, 10.8939, 7.205796, 
    2.473217,
  -0.6725413, -2.512176, -5.647513, -10.26797, -15.63438, -20.13788, 
    -21.51631, -18.58341, -12.98447, -7.37911, -3.116992, -2.430194e-05, 
    3.11676, 7.377151, 12.97045, 18.50855, 21.20838, 19.1347, 12.99875, 
    4.582281,
  -1.864758, -6.489053, -13.15883, -21.46106, -29.61354, -35.64208, 
    -37.64965, -33.83036, -25.30485, -15.61154, -7.108466, -7.180536e-05, 
    7.107486, 15.60288, 25.24927, 33.56337, 36.65423, 32.71277, 22.70754, 
    8.173388,
  -4.30142, -14.02004, -25.7063, -37.56685, -46.92198, -52.71651, -55.25098, 
    -51.81897, -41.29388, -27.32007, -13.2053, -0.0002546461, 13.2018, 
    27.29113, 41.12322, 51.05972, 52.63205, 45.65824, 31.83648, 11.54705,
  -8.382675, -25.65773, -42.53046, -55.63113, -63.05907, -66.50754, 
    -69.94808, -69.17681, -58.78362, -41.37749, -20.97836, -0.0007577671, 
    20.96911, 41.30459, 58.37036, 67.41364, 64.20592, 52.21219, 35.23764, 
    12.525,
  -14.264, -41.12642, -61.88537, -73.0153, -76.14981, -76.48225, -81.86056, 
    -86.18807, -78.16755, -58.14941, -30.63301, -0.001274176, 30.61667, 
    58.01537, 77.37727, 82.75978, 71.04005, 51.32878, 31.31981, 10.27485,
  -24.23621, -68.90245, -101.6995, -118.0156, -120.1859, -113.4333, 
    -106.7686, -97.85954, -80.78855, -56.91515, -29.1768, -0.000617792, 
    29.16827, 56.8361, 80.23028, 94.73743, 92.57227, 74.5586, 48.76833, 
    16.5039,
  -31.92004, -89.28856, -128.6348, -146.5004, -149.2513, -145.0696, 
    -140.8036, -130.0807, -107.3828, -75.52354, -38.7186, -0.0006360901, 
    38.70978, 75.44006, 106.7683, 126.4058, 122.8486, 94.79347, 57.64728, 
    18.50382,
  -37.62951, -104.9204, -150.4181, -170.9715, -175.5504, -174.9853, 
    -171.2431, -155.8773, -127.5584, -89.47076, -45.9027, -0.0007478549, 
    45.89281, 89.38064, 126.9091, 151.9632, 151.0847, 116.7305, 68.70924, 
    21.58605,
  -41.16886, -115.0286, -165.3458, -188.5078, -194.612, -196.2929, -192.0633, 
    -173.1506, -141.1849, -99.028, -50.87502, -0.0008732486, 50.86376, 
    98.9285, 140.4886, 169.0364, 170.6394, 133.2431, 77.92146, 24.42149,
  -42.92503, -120.316, -173.7073, -198.8369, -205.9526, -208.4872, -203.7117, 
    -183.0177, -149.1435, -104.6862, -53.83649, -0.0009701027, 53.82409, 
    104.5784, 148.4046, 178.7401, 181.6155, 143.0701, 84.05826, 26.47159,
  -43.4308, -121.9028, -176.3468, -202.2156, -209.6905, -212.391, -207.4106, 
    -186.2277, -151.7736, -106.5698, -54.82485, -0.001038348, 54.81197, 
    106.4588, 151.0177, 181.8859, 185.1004, 146.2845, 86.21567, 27.22481,
  -42.92503, -120.316, -173.7075, -198.8372, -205.9531, -208.4873, -203.7117, 
    -183.0177, -149.1436, -104.6863, -53.83656, -0.0009746035, 53.82415, 
    104.5786, 148.4047, 178.7402, 181.6154, 143.0701, 84.05879, 26.47186,
  -41.16894, -115.0291, -165.3479, -188.513, -194.6198, -196.2951, -192.0631, 
    -173.1521, -141.1867, -99.02976, -50.87612, -0.0008743054, 50.86488, 
    98.93025, 140.4904, 169.0376, 170.6385, 133.2451, 77.92902, 24.42477,
  -37.63055, -104.9261, -150.4367, -171.0152, -175.6185, -175.0226, 
    -171.2572, -155.8947, -127.5757, -89.48642, -45.91221, -0.0007228057, 
    45.90232, 89.39616, 126.9259, 151.9783, 151.0945, 116.7676, 68.77449, 
    21.61243,
  -31.92789, -89.32772, -128.7533, -146.7651, -149.6796, -145.4587, 
    -141.0587, -130.2592, -107.5229, -75.63213, -38.78001, -0.0006301514, 
    38.7711, 75.54806, 106.905, 126.5723, 123.0885, 95.1803, 58.04871, 
    18.65579,
  -24.27981, -69.10388, -102.2662, -119.2233, -122.1702, -115.8263, 
    -108.7934, -99.24502, -81.75626, -57.54005, -29.48654, -0.0006429676, 
    29.47774, 57.45884, 81.18667, 96.09075, 94.56637, 76.91576, 50.58172, 
    17.15991,
  -14.44595, -41.90964, -63.93599, -77.18231, -82.96422, -85.58506, 
    -91.41525, -94.00819, -83.45747, -61.19652, -31.98156, -0.001369348, 
    31.96444, 61.05779, 82.64923, 90.53899, 80.51928, 60.20017, 37.35996, 
    12.39852,
  -8.991517, -28.10656, -48.46344, -66.88348, -80.4401, -88.95592, -94.00536, 
    -90.06506, -73.66981, -50.18956, -24.88999, -0.0008415745, 24.87985, 
    50.11125, 73.23431, 88.22974, 88.01983, 73.8138, 50.10574, 17.82771,
  -5.957871, -20.21561, -39.39774, -61.36924, -81.04043, -94.73871, 
    -100.3594, -92.57339, -71.76904, -46.09989, -21.74741, -0.0003320602, 
    21.7432, 46.06514, 71.56295, 91.6395, 97.01472, 85.24337, 59.46204, 
    21.55882,
  -0.9399071, -3.336047, -7.072988, -12.34265, -18.40515, -23.57117, 
    -25.37567, -22.44798, -16.34557, -9.797296, -4.360099, -0.0001434187, 
    4.358913, 9.789782, 16.30696, 22.28852, 24.83702, 22.05953, 14.84148, 
    5.202405,
  -1.981441, -6.567601, -12.58139, -19.77936, -26.96574, -32.5401, -34.56007, 
    -31.46413, -24.24913, -15.62514, -7.43037, -0.00060021, 7.42574, 
    15.59845, 24.12655, 31.01145, 33.19006, 29.10857, 19.78053, 7.013086,
  -4.235604, -13.26424, -23.20453, -32.99271, -41.07483, -46.56984, -48.9064, 
    -46.01409, -37.43953, -25.64855, -12.83404, -0.002207298, 12.81828, 
    25.56509, 37.08536, 44.80064, 45.5069, 38.76159, 26.23974, 9.319622,
  -7.867774, -23.41737, -37.69667, -48.87862, -56.11146, -60.28139, 
    -63.11863, -61.63081, -52.67139, -37.87604, -19.66004, -0.006301285, 
    19.61759, 37.66442, 51.8212, 58.87393, 55.87303, 44.89161, 29.36364, 
    10.21294,
  -12.70405, -36.05611, -53.69087, -63.97278, -68.42944, -70.36257, -74.2143, 
    -75.76202, -68.0305, -51.05072, -27.27573, -0.01382015, 27.18572, 
    50.61371, 66.31303, 70.36181, 60.74961, 43.85423, 26.24308, 8.551584,
  -18.37201, -49.9237, -69.32902, -76.852, -77.77195, -77.49903, -83.12653, 
    -89.31077, -84.44051, -65.97806, -36.14514, -0.02120624, 36.00262, 
    65.2563, 81.49487, 79.95569, 60.685, 36.39178, 17.68551, 4.725903,
  -28.35539, -76.36891, -105.0195, -115.4847, -114.3165, -106.7582, 
    -100.7411, -95.08454, -82.43252, -61.29976, -32.77573, -0.01015503, 
    32.7011, 60.86786, 80.31308, 86.53587, 72.84867, 48.21571, 26.39515, 
    7.845399,
  -36.01314, -95.69952, -129.2956, -140.7802, -140.419, -135.2433, -131.7582, 
    -125.8042, -108.927, -80.41544, -42.74271, -0.009889354, 42.6684, 
    79.96743, 106.5816, 115.572, 96.61889, 60.95701, 30.35975, 8.314462,
  -42.55059, -112.4489, -150.9757, -164.258, -165.6228, -164.0838, -161.8129, 
    -152.2676, -130.0041, -95.05602, -50.27802, -0.01091109, 50.19876, 
    94.58942, 127.5634, 141.2508, 121.7647, 77.24188, 36.94234, 9.794385,
  -47.38434, -125.0041, -167.5573, -182.4497, -185.1595, -186.5025, 
    -184.2627, -171.0429, -144.7459, -105.3275, -55.59187, -0.01240995, 
    55.50434, 104.8271, 142.1834, 159.496, 141.107, 90.92146, 42.82894, 
    11.23961,
  -50.28202, -132.6694, -177.9348, -194.0039, -197.5119, -200.4399, 
    -197.8248, -182.243, -153.6114, -111.57, -58.84203, -0.01373562, 
    58.74681, 111.0362, 150.9283, 170.3048, 152.9473, 99.88643, 46.98642, 
    12.34098,
  -51.2363, -135.2286, -181.4612, -197.9704, -201.7394, -205.1441, -202.342, 
    -185.979, -156.5931, -113.6835, -59.94629, -0.01430562, 59.84787, 
    113.1357, 153.8596, 173.8899, 156.9101, 102.9979, 48.49813, 12.75777,
  -50.2823, -132.6707, -177.9385, -194.0111, -197.5205, -200.4404, -197.823, 
    -182.244, -153.6132, -111.5718, -58.8432, -0.01376611, 58.74794, 
    111.0379, 150.9298, 170.3051, 152.9439, 99.88657, 46.99446, 12.34491,
  -47.38671, -125.0143, -167.5834, -182.499, -185.2215, -186.52, -184.2608, 
    -171.0527, -144.7588, -105.3403, -55.59998, -0.01240825, 55.5124, 
    104.8396, 142.1945, 159.5005, 141.0964, 90.93815, 42.88594, 11.26535,
  -42.56501, -112.5074, -151.1174, -164.5192, -165.9705, -164.284, -161.8992, 
    -152.3555, -130.0882, -95.1313, -50.32384, -0.01091776, 50.24423, 
    94.66243, 127.6378, 141.3124, 121.8203, 77.44056, 37.25428, 9.924028,
  -36.08174, -95.96466, -129.9068, -141.8836, -141.9692, -136.6675, -132.768, 
    -126.514, -109.4656, -80.81993, -42.96814, -0.01013835, 42.89202, 
    80.36219, 107.0826, 116.1996, 97.56167, 62.34772, 31.70666, 8.833057,
  -28.61595, -77.33565, -107.143, -119.2032, -119.6793, -113.0126, -106.2635, 
    -99.131, -85.38991, -63.25858, -33.75848, -0.01094862, 33.67863, 
    62.80209, 83.18985, 90.43469, 78.24883, 54.19913, 30.88222, 9.485172,
  -19.16233, -52.74026, -75.2159, -86.77852, -91.99849, -95.2523, -101.864, 
    -105.68, -96.60992, -73.6897, -39.81519, -0.02319499, 39.66205, 72.92961, 
    93.56616, 96.13721, 79.01505, 52.9949, 29.01985, 8.752895,
  -14.71346, -42.92911, -67.23377, -85.42661, -97.49469, -105.2572, 
    -111.4269, -109.8444, -94.63405, -68.58049, -35.81927, -0.01603512, 
    35.71755, 68.09961, 92.78214, 104.0591, 96.80927, 75.56881, 48.01914, 
    16.34579,
  -12.14072, -37.35803, -63.31583, -86.576, -103.9607, -115.3617, -121.8546, 
    -117.2139, -97.9218, -68.90224, -35.21702, -0.008146606, 35.16262, 
    68.63239, 96.82998, 113.5794, 111.8377, 92.78121, 62.08585, 21.93482,
  -2.585937, -8.402172, -15.72178, -24.3613, -33.10421, -40.12339, -43.00172, 
    -39.82972, -31.54926, -20.98549, -10.25333, -0.002723871, 10.23773, 
    20.91673, 31.29331, 39.03057, 40.88101, 35.30836, 23.69003, 8.334777,
  -4.197906, -12.96253, -22.38141, -31.83899, -40.21106, -46.39047, 
    -48.99966, -46.10712, -37.76741, -26.19143, -13.26731, -0.008377265, 
    13.22358, 26.01703, 37.17415, 44.41043, 44.8836, 37.89876, 25.21059, 
    8.839775,
  -7.183688, -21.17375, -33.82354, -44.06836, -51.44724, -56.24746, 
    -58.80894, -56.79446, -48.4463, -35.06224, -18.35453, -0.02320621, 
    18.241, 34.63832, 47.08615, 53.132, 50.51359, 40.47753, 26.06722, 8.967216,
  -11.09512, -31.47951, -47.17439, -57.21511, -62.73808, -65.80451, 
    -68.79256, -68.57649, -60.77049, -45.4993, -24.37728, -0.05300032, 
    24.12894, 44.6115, 58.03048, 61.52069, 53.72737, 39.24822, 23.48246, 
    7.680413,
  -15.22176, -41.85984, -59.57104, -68.29033, -71.43699, -72.7384, -76.67151, 
    -79.26414, -72.96049, -56.29274, -30.72708, -0.09832585, 30.27386, 
    54.69427, 68.09404, 67.07327, 51.98256, 32.36716, 16.53432, 4.744534,
  -19.00507, -51.00944, -69.79496, -76.81236, -77.86185, -77.80381, 
    -83.21006, -89.57743, -85.84931, -68.27873, -37.93253, -0.1397676, 
    37.26662, 65.82668, 78.13761, 70.24601, 45.83812, 21.07819, 6.660569, 
    0.8250513,
  -26.95016, -72.40556, -99.3354, -109.1824, -108.1344, -100.9968, -95.23047, 
    -90.72768, -80.27201, -61.04369, -33.16236, -0.0681086, 32.80616, 
    59.53056, 74.56389, 72.96306, 51.02629, 25.82205, 10.90776, 2.564681,
  -32.58745, -87.13342, -118.9035, -130.8113, -131.353, -126.5672, -123.0984, 
    -118.995, -105.4035, -79.52568, -42.86052, -0.06423534, 42.51222, 
    77.95262, 98.96931, 97.40909, 68.04713, 33.57568, 12.77789, 2.653711,
  -37.94156, -101.1902, -137.7678, -152.0002, -154.7408, -153.6081, 
    -151.6815, -144.8783, -126.2578, -93.91965, -50.18457, -0.06708392, 
    49.82836, 92.32221, 119.5699, 121.2392, 88.38724, 44.99184, 16.7554, 
    3.435803,
  -42.39817, -112.8185, -153.2132, -169.1594, -173.6395, -175.9124, 
    -174.4707, -164.0875, -141.1107, -104.009, -55.29734, -0.07326273, 
    54.91868, 102.351, 134.2143, 139.2337, 105.4783, 55.24656, 20.26129, 
    4.105556,
  -45.39536, -120.6042, -163.4821, -180.4691, -186.0044, -190.5122, 
    -188.9369, -175.8249, -150.0868, -110.1171, -58.40384, -0.07928593, 
    58.00132, 108.3882, 142.988, 150.2248, 116.6354, 62.34725, 22.72892, 
    4.58338,
  -46.45689, -123.3563, -167.1013, -184.4393, -190.3228, -195.5841, 
    -193.8788, -179.7787, -153.1083, -112.1808, -59.45667, -0.08181569, 
    59.04398, 110.4208, 145.9225, 153.9118, 120.4907, 64.88472, 23.63068, 
    4.761972,
  -45.39927, -120.6185, -163.5124, -180.5173, -186.0545, -190.5148, 
    -188.9253, -175.8286, -150.0947, -110.1258, -58.40948, -0.07934053, 
    58.00672, 108.3959, 142.9925, 150.2196, 116.6113, 62.34824, 22.77194, 
    4.604698,
  -42.41886, -112.8914, -153.363, -169.3955, -173.9019, -175.9932, -174.4681, 
    -164.1228, -141.1558, -104.0542, -55.32612, -0.07347433, 54.94623, 
    102.3909, 134.241, 139.2274, 105.4312, 55.32468, 20.48188, 4.205576,
  -38.02903, -101.4902, -138.365, -152.9384, -155.8632, -154.3035, -152.0321, 
    -145.1797, -126.5157, -94.1377, -50.31483, -0.06810629, 49.95296, 
    92.51685, 119.7543, 121.4048, 88.6306, 45.66079, 17.66846, 3.814526,
  -32.89396, -88.15829, -120.8846, -133.9034, -135.3034, -130.2738, 
    -125.9313, -121.0352, -106.899, -80.5864, -43.43187, -0.06813898, 
    43.06387, 78.93997, 100.2681, 99.16269, 70.68756, 37.02671, 15.85981, 
    3.833008,
  -27.84833, -75.33356, -104.8026, -117.5323, -119.1202, -113.5009, 
    -106.6412, -99.57543, -86.98579, -65.57291, -35.45167, -0.07733482, 
    35.05381, 63.92685, 80.97136, 81.4006, 62.00542, 37.12965, 19.04383, 
    5.510602,
  -21.17696, -57.90607, -82.18564, -95.12104, -101.7338, -106.1548, 
    -113.1733, -116.8768, -107.4252, -82.80888, -45.16869, -0.1573081, 
    44.43742, 80.19238, 99.37449, 96.88381, 74.23958, 45.69691, 23.05624, 
    6.587244,
  -19.74832, -55.81491, -83.41969, -101.5452, -112.5475, -119.6886, 
    -126.4634, -126.3286, -111.7281, -83.39633, -44.57574, -0.1173594, 
    44.05037, 81.59702, 106.33, 112.7265, 98.0842, 70.98228, 42.08015, 
    13.68623,
  -19.11134, -55.39455, -85.8554, -107.8918, -122.0605, -131.2246, -138.1727, 
    -135.9726, -118.2829, -87.09834, -46.15498, -0.0719446, 45.82209, 
    85.9129, 114.5687, 126.0403, 115.6982, 88.9489, 55.43679, 18.65927,
  -7.048122, -21.22888, -35.31716, -48.50101, -59.73624, -68.09098, 
    -72.09499, -69.20831, -58.72572, -42.36473, -22.14648, -0.06409311, 
    21.90062, 41.64902, 56.81775, 64.74842, 62.93559, 51.58811, 33.57413, 
    11.6319,
  -8.535301, -25.00342, -39.75827, -52.01344, -61.48125, -68.10502, 
    -71.36241, -68.76495, -58.88569, -42.92951, -22.64144, -0.1311353, 
    22.16844, 41.65269, 55.70341, 61.82053, 58.11279, 46.03846, 29.18475, 
    9.942898,
  -10.83522, -30.84708, -46.72679, -57.83725, -65.03993, -69.50156, 
    -72.20586, -70.52205, -61.56522, -45.72751, -24.46459, -0.2657216, 
    23.54097, 43.35048, 55.90898, 58.83554, 51.3862, 37.57775, 22.35461, 
    7.301213,
  -13.00739, -36.38531, -53.43458, -63.72355, -69.16184, -71.9427, -74.72463, 
    -74.58541, -66.72174, -50.58696, -27.46234, -0.4801658, 25.82883, 
    46.49828, 57.27399, 55.85566, 43.305, 27.31181, 14.24638, 4.21325,
  -14.29367, -39.75961, -57.72796, -67.76132, -72.29939, -74.10948, 
    -77.49841, -79.36996, -72.89937, -56.42882, -31.06225, -0.7571421, 
    28.49436, 50.02781, 58.27302, 51.23397, 32.86592, 15.22503, 5.298873, 
    0.925532,
  -14.45004, -40.44544, -59.17139, -69.78371, -74.50197, -76.11981, 
    -80.50135, -84.70364, -79.98994, -63.27407, -35.2995, -1.003393, 
    31.78786, 54.16396, 58.756, 44.47916, 20.13189, 2.142166, -3.65747, 
    -2.215316,
  -18.59665, -52.77212, -78.44942, -92.71613, -96.28255, -91.93681, 
    -86.54606, -81.35529, -71.35331, -54.15801, -29.52128, -0.511152, 
    27.55172, 48.20391, 54.93338, 44.34748, 19.88392, 2.533029, -1.821058, 
    -1.184787,
  -20.53482, -59.02592, -89.42015, -107.8729, -114.7321, -113.1519, -109.568, 
    -104.7514, -92.68892, -70.2649, -38.07952, -0.4754617, 36.14543, 
    63.89416, 73.5575, 59.46222, 29.01142, 7.344388, -0.1036701, -0.7921886,
  -22.7091, -65.84892, -101.0246, -123.6467, -134.1196, -136.3556, -134.3759, 
    -127.8015, -111.6662, -83.41063, -44.7155, -0.4659536, 42.81808, 
    77.00503, 91.37955, 77.05575, 41.9029, 14.69072, 2.761814, -0.08894855,
  -24.69319, -71.91061, -110.9898, -136.888, -150.4404, -156.5509, -155.5387, 
    -146.0267, -125.6445, -92.62803, -49.25649, -0.4759242, 47.34988, 
    86.22444, 104.8911, 91.98138, 53.88393, 21.39535, 5.035598, 0.3792426,
  -26.13708, -76.23483, -117.9147, -145.9156, -161.5266, -170.4274, 
    -169.6807, -157.5284, -134.1149, -98.09869, -51.93346, -0.4923958, 
    49.98998, 91.64943, 113.1177, 101.7309, 62.31421, 26.19577, 6.589716, 
    0.6762621,
  -26.6794, -77.84406, -120.4609, -149.2019, -165.5263, -175.371, -174.6124, 
    -161.44, -136.9534, -99.92392, -52.8273, -0.5003834, 50.86335, 93.44178, 
    115.8563, 105.0701, 65.29958, 27.93827, 7.189875, 0.8018587,
  -26.18473, -76.3828, -118.1679, -146.2472, -161.8276, -170.4534, -169.6116, 
    -157.5306, -134.1375, -98.12825, -51.95423, -0.4941755, 50.00344, 
    91.65562, 113.08, 101.6363, 62.16683, 26.21022, 6.801472, 0.7807001,
  -24.86576, -72.44231, -111.894, -138.0898, -151.6322, -157.0078, -155.6122, 
    -146.1676, -125.7823, -92.75871, -49.34132, -0.4835996, 47.40372, 
    86.26141, 104.8124, 91.83447, 53.76776, 21.78304, 5.854045, 0.745253,
  -23.22259, -67.41748, -103.673, -127.2188, -137.9963, -139.0749, -136.0568, 
    -129.0645, -112.5614, -84.05007, -45.07471, -0.4926394, 43.07507, 
    77.36608, 91.72881, 77.73831, 43.20846, 16.96348, 5.317594, 0.9493166,
  -21.85169, -63.00449, -96.05582, -116.8835, -125.2396, -123.3367, 
    -118.0502, -111.1815, -97.35594, -73.36204, -39.66904, -0.5433602, 
    37.49714, 66.43572, 77.31298, 65.04762, 36.6128, 15.59244, 6.456908, 
    1.657174,
  -21.51344, -61.44365, -92.58012, -111.6635, -119.0184, -117.0832, 
    -110.1774, -100.7411, -86.68986, -64.77978, -34.97682, -0.6200627, 
    32.66644, 58.13577, 69.18432, 62.43684, 41.19972, 22.19052, 11.31303, 
    3.430954,
  -19.91998, -56.41972, -84.49461, -102.9197, -113.9427, -120.6815, 
    -127.3692, -128.7366, -116.4812, -89.03004, -48.59534, -1.158748, 
    44.65883, 79.15189, 93.78325, 85.3699, 60.22007, 34.1786, 16.30948, 
    4.543395,
  -23.36438, -65.64289, -97.15734, -117.0361, -128.5127, -135.4804, 
    -141.8534, -141.2203, -125.5486, -94.53384, -51.06623, -0.9285723, 
    47.99419, 87.0359, 108.3447, 107.0868, 84.6252, 54.51537, 28.98041, 
    8.739227,
  -25.99702, -72.65333, -106.6677, -127.5178, -139.3536, -146.6876, 
    -153.0588, -151.3371, -133.6431, -100.1131, -53.85308, -0.6797881, 
    51.55476, 94.31158, 119.786, 122.3226, 101.0085, 67.90187, 37.02478, 
    11.32684,
  -10.76042, -31.52585, -50.12208, -65.52389, -77.37614, -85.69749, 
    -89.78414, -86.76494, -74.89243, -55.11389, -29.3095, -0.2934685, 
    28.36186, 52.87218, 69.81956, 76.48459, 71.23688, 56.05466, 35.30945, 
    11.9933,
  -11.30003, -32.67904, -50.86678, -64.98934, -75.21021, -81.99158, 
    -85.30885, -82.43174, -71.22584, -52.48618, -27.99371, -0.4990779, 
    26.4544, 49.074, 63.95594, 68.59418, 61.96783, 47.19435, 29.00336, 
    9.697211,
  -11.98483, -34.21598, -52.07566, -64.7724, -73.02286, -77.86364, -80.47907, 
    -78.26582, -68.17719, -50.62656, -27.24061, -0.8738182, 24.61977, 
    45.06352, 56.86259, 57.92404, 48.53173, 34.0298, 19.644, 6.299206,
  -12.19171, -34.72129, -52.49216, -64.51736, -71.59516, -75.0698, -77.53415, 
    -76.50915, -67.70941, -50.98505, -27.81615, -1.416038, 23.62797, 
    42.30038, 50.56232, 47.01657, 34.0628, 19.9115, 9.8435, 2.796536,
  -11.51238, -33.16, -50.87915, -63.16758, -70.23205, -73.25797, -76.13326, 
    -76.62816, -69.23037, -53.06065, -29.41628, -2.072119, 23.28211, 40.3658, 
    44.50259, 35.52853, 18.98224, 5.897589, 0.5706131, -0.4229418,
  -9.900175, -29.36697, -46.97984, -60.49796, -68.82292, -72.40363, 
    -76.09712, -78.16738, -72.17252, -56.34908, -31.69348, -2.664317, 
    23.58012, 38.95861, 37.95737, 22.71407, 3.40764, -7.239598, -7.53751, 
    -3.113432,
  -12.23918, -36.8522, -59.85234, -76.92087, -84.80756, -83.71325, -79.26623, 
    -73.20171, -62.79891, -46.97913, -25.65408, -1.408306, 20.93523, 
    35.17458, 35.73478, 22.52571, 2.363383, -7.407221, -6.170084, -2.271746,
  -12.50472, -38.70692, -65.35012, -87.14435, -99.33399, -101.5426, 
    -98.81557, -92.92136, -80.92454, -60.91942, -33.15083, -1.321714, 
    28.43853, 47.9629, 48.89062, 31.34594, 8.270387, -2.875101, -3.854155, 
    -1.546273,
  -13.03403, -41.23544, -71.7076, -98.31039, -115.0732, -121.368, -120.3425, 
    -113.231, -98.01846, -72.99343, -39.29027, -1.261746, 34.7154, 59.82275, 
    63.39643, 43.70135, 17.42165, 3.412739, -0.8025614, -0.6371123,
  -13.53034, -43.48449, -77.18626, -107.8383, -128.6475, -139.0402, 
    -139.3348, -130.0526, -111.1507, -81.68631, -43.54725, -1.239273, 
    39.07729, 68.63901, 75.46092, 55.33173, 26.29742, 8.984547, 1.566632, 
    -0.0008243099,
  -13.91593, -45.14609, -81.09354, -114.5175, -138.1316, -151.4889, 
    -152.3981, -140.9829, -119.233, -86.8377, -46.02755, -1.243856, 41.58496, 
    73.8912, 83.1694, 63.44837, 32.78406, 12.97616, 3.196094, 0.4219927,
  -14.09409, -45.85816, -82.67225, -117.117, -141.7019, -155.9822, -156.9837, 
    -144.7288, -121.9414, -88.5443, -46.84822, -1.251653, 42.39658, 75.60267, 
    85.73858, 66.25694, 35.06043, 14.41886, 3.870849, 0.6184167,
  -14.06136, -45.57763, -81.77905, -115.3478, -138.8467, -151.5925, 
    -152.2558, -140.962, -119.2451, -86.86906, -46.05598, -1.255983, 
    41.56948, 73.80753, 82.95586, 63.17186, 32.48483, 13.01871, 3.610784, 
    0.6251337,
  -13.97877, -44.81362, -79.3049, -110.4657, -131.1429, -140.1693, -139.6652, 
    -130.3712, -111.3732, -81.865, -43.66882, -1.284828, 39.04079, 68.44009, 
    75.0412, 55.0476, 26.26404, 9.770172, 2.984144, 0.6251461,
  -14.16217, -44.56961, -77.02843, -105.0601, -122.1284, -126.7101, 
    -123.9941, -115.9184, -99.80669, -74.13032, -39.90102, -1.391946, 
    34.90701, 60.09286, 63.95478, 45.40595, 20.20433, 7.222829, 3.042779, 
    0.8970752,
  -14.97276, -45.95362, -76.85246, -101.9293, -115.9387, -117.9046, -112.958, 
    -103.9776, -89.09204, -66.28851, -35.89221, -1.58369, 30.42028, 52.0062, 
    55.4114, 40.94662, 20.06444, 8.631376, 4.671801, 1.567624,
  -16.93861, -50.48471, -81.13422, -104.1099, -116.2096, -117.9129, 
    -111.6922, -100.3684, -84.66841, -62.36174, -33.68153, -1.747245, 
    28.0667, 49.12832, 55.61877, 46.94391, 29.27937, 15.76576, 8.480619, 
    2.737551,
  -17.52581, -51.2179, -80.47507, -102.664, -117.3784, -126.0961, -132.1766, 
    -131.1686, -116.665, -88.20736, -48.38583, -3.09732, 39.20039, 69.0541, 
    79.03157, 68.54653, 45.88356, 24.77379, 11.34772, 3.065735,
  -22.55229, -64.24941, -97.15991, -119.5002, -133.0302, -140.6732, 
    -146.0817, -143.6235, -126.3943, -94.6293, -51.40986, -2.574466, 
    43.90643, 79.2204, 95.76529, 90.26762, 66.68555, 39.49694, 19.35557, 
    5.474343,
  -26.07633, -73.29076, -108.6111, -131.0959, -144.0987, -151.3958, 
    -156.5166, -153.0989, -134.0654, -99.92576, -53.95684, -2.041567, 
    47.89873, 87.08158, 107.538, 104.6112, 80.22693, 49.0351, 24.35888, 
    6.934532,
  -15.28871, -44.02893, -68.00451, -86.00657, -98.41114, -106.0656, 
    -109.1042, -104.5566, -90.0755, -66.44455, -35.78997, -1.65509, 31.29922, 
    58.13554, 74.67024, 78.3319, 68.84061, 50.76294, 30.23171, 9.906862,
  -13.97598, -40.42244, -62.84236, -79.93329, -91.67974, -98.60754, 
    -101.2468, -96.95464, -83.38723, -61.47506, -33.33879, -2.330028, 
    27.21552, 50.7575, 64.58131, 66.68581, 57.35574, 41.52874, 24.57408, 
    8.02677,
  -11.94078, -34.89123, -55.06604, -70.96006, -81.89265, -87.8765, -90.17936, 
    -86.61474, -74.60136, -55.15655, -30.3752, -3.466761, 21.46805, 40.24348, 
    49.76561, 49.05193, 39.52606, 26.9489, 15.51687, 4.980974,
  -9.497222, -28.35352, -46.17593, -61.1904, -71.78047, -77.21261, -79.52341, 
    -77.04832, -66.84206, -49.86675, -28.16373, -4.978326, 15.50863, 
    29.19958, 33.667, 29.4345, 19.61852, 10.80018, 5.537479, 1.629369,
  -6.769984, -21.10356, -36.55006, -51.17192, -62.23327, -67.958, -70.75489, 
    -69.52783, -61.12924, -46.30898, -27.00795, -6.709813, 9.924904, 
    18.54064, 17.49352, 9.50826, -0.1036429, -4.646647, -3.800922, -1.464018,
  -3.783877, -13.1788, -26.22869, -41.0714, -53.68618, -60.81796, -64.5021, 
    -64.31246, -57.38709, -44.1943, -26.55323, -8.358675, 4.82612, 8.037785, 
    0.8735638, -10.52252, -18.34259, -17.7116, -11.29999, -3.857783,
  -4.630501, -15.96399, -31.31317, -47.97113, -60.46613, -65.21684, 
    -64.22437, -58.31573, -48.06508, -35.00824, -19.84727, -4.7036, 6.494187, 
    9.311674, 2.560287, -8.681206, -18.13177, -17.45971, -10.26803, -3.251176,
  -3.756479, -14.15864, -30.70683, -50.86903, -67.8858, -76.55929, -77.7538, 
    -72.20221, -60.96798, -45.1953, -25.40514, -4.558962, 11.59389, 16.05541, 
    6.751253, -7.204104, -14.91313, -12.95262, -7.30093, -2.202868,
  -3.144104, -13.07473, -31.14913, -55.05592, -76.87529, -89.98496, 
    -93.53105, -87.82042, -74.73534, -55.41272, -30.71095, -4.301955, 
    17.17794, 24.87399, 14.77912, -1.697031, -9.22126, -7.372427, -3.886547, 
    -1.041388,
  -2.610243, -12.13187, -31.5601, -58.82092, -85.04196, -102.4353, -108.1772, 
    -101.8681, -86.41628, -63.51697, -34.71466, -4.064769, 21.72275, 
    32.91646, 23.35628, 4.891892, -3.573169, -2.671859, -1.199888, -0.1596564,
  -2.295743, -11.64834, -32.13421, -61.82887, -91.173, -111.5593, -118.6886, 
    -111.5461, -94.00722, -68.50022, -37.0981, -3.93499, 24.48592, 38.20691, 
    29.61849, 10.1006, 0.6482382, 0.6166029, 0.6782439, 0.4574451,
  -2.307762, -11.83673, -32.89093, -63.54084, -93.8991, -114.9615, -122.3632, 
    -114.8891, -96.55013, -70.13152, -37.87841, -3.923049, 25.31175, 
    39.83266, 31.61625, 11.82697, 1.987043, 1.755352, 1.519073, 0.767122,
  -2.762821, -12.99265, -34.15832, -64.13675, -93.11095, -112.1197, 
    -118.5014, -111.4435, -93.90072, -68.43948, -37.11098, -4.057119, 
    24.1334, 37.48438, 28.71708, 9.462959, 0.1292934, 0.695713, 1.400326, 
    0.810178,
  -3.819301, -15.6199, -36.86178, -65.05054, -90.82285, -105.7591, -109.7086, 
    -102.8936, -86.91766, -63.75497, -34.92245, -4.432704, 20.90683, 
    31.54113, 22.19121, 4.864069, -3.093692, -1.239421, 0.9738659, 0.7821808,
  -5.627882, -20.24892, -42.14157, -68.36541, -90.46497, -101.3242, 
    -102.1359, -94.24958, -79.07634, -58.02937, -32.15601, -5.07367, 
    16.68011, 24.90995, 16.73876, 2.863594, -3.741078, -1.652668, 1.114561, 
    0.8882958,
  -8.181149, -26.92606, -50.34206, -75.17447, -94.47768, -103.2799, 
    -101.6614, -91.51617, -75.7849, -55.21246, -30.76699, -5.670527, 
    14.40593, 23.05747, 18.50141, 8.272887, 1.473753, 1.016668, 1.982992, 
    1.043396,
  -11.48754, -35.6708, -61.52, -85.62222, -102.918, -110.8264, -107.7525, 
    -95.39009, -78.33525, -56.73173, -31.57951, -5.837038, 15.68198, 
    27.75553, 28.13655, 20.59394, 11.26142, 5.52334, 2.917695, 1.016641,
  -12.82959, -39.19137, -66.1949, -91.17905, -110.7379, -122.9218, -128.6268, 
    -124.8006, -108.4473, -81.19177, -46.43201, -9.77728, 21.33699, 39.64614, 
    41.84076, 31.7028, 17.51299, 6.945755, 1.875549, 0.1751231,
  -17.42289, -51.66493, -83.23718, -109.1236, -127.2159, -137.1902, 
    -141.4222, -136.1257, -117.3727, -87.13012, -49.02254, -8.540474, 
    27.2267, 51.01121, 58.11761, 49.37118, 31.00403, 14.40143, 5.253628, 
    1.04487,
  -20.24779, -59.4005, -94.01149, -120.8752, -138.5825, -147.587, -150.849, 
    -144.2404, -123.5864, -91.11271, -50.56955, -7.388656, 31.44061, 
    58.48723, 68.25933, 60.2207, 39.73294, 19.76616, 7.944012, 1.820552,
  -16.37654, -47.28059, -73.27827, -92.84277, -105.9676, -113.2491, 
    -115.1323, -109.0247, -92.96806, -68.27567, -37.4164, -4.028646, 
    27.32307, 51.91567, 65.93414, 67.45426, 57.06767, 40.27166, 23.13363, 
    7.403176,
  -14.32957, -41.75707, -65.66742, -84.40087, -97.28205, -104.3419, 
    -106.2815, -100.8191, -86.02687, -63.35376, -35.25349, -5.192288, 
    22.58197, 43.82912, 55.39222, 56.03564, 46.70488, 32.70493, 18.92619, 
    6.092268,
  -11.21575, -33.29695, -53.89785, -71.26786, -83.79737, -90.61651, 
    -92.83655, -88.60608, -75.89222, -56.29473, -32.26425, -7.10032, 
    15.30884, 31.36504, 38.90301, 37.83533, 29.80871, 20.02366, 11.62488, 
    3.749725,
  -7.754339, -23.81077, -40.55894, -56.33614, -68.61984, -75.45789, 
    -78.20534, -75.49262, -65.19653, -49.0107, -29.39169, -9.572368, 
    6.803576, 16.77959, 19.41649, 16.19617, 9.748762, 4.924914, 2.77684, 
    0.8686572,
  -4.300157, -14.24601, -26.95358, -41.11857, -53.49488, -60.95619, 
    -64.51161, -63.2832, -55.37174, -42.46559, -27.02712, -12.37702, 
    -2.147658, 1.279613, -1.465755, -6.780653, -10.92164, -10.26956, 
    -6.137635, -2.035426,
  -0.9411106, -4.888021, -13.61916, -26.47457, -39.64539, -48.65001, 
    -53.24036, -53.08695, -47.11676, -36.93845, -25.08334, -15.18881, 
    -11.21653, -14.94396, -23.33582, -29.81977, -29.91165, -23.15666, 
    -13.46165, -4.363004,
  -1.272845, -5.807214, -14.95761, -27.91246, -40.47945, -48.38496, 
    -50.90304, -46.88976, -38.04528, -27.60919, -17.19083, -8.942434, 
    -5.897779, -9.981384, -18.68163, -25.86241, -28.17102, -22.37177, 
    -12.60141, -3.911275,
  -0.2196815, -3.101723, -12.01797, -26.82627, -42.89134, -54.4634, 
    -59.63766, -56.61874, -47.31234, -35.04417, -21.25871, -8.932316, 
    -3.211668, -8.103115, -19.78158, -27.58084, -26.21497, -18.3661, 
    -9.715528, -2.859698,
  0.511555, -1.30722, -10.43316, -27.38816, -47.22294, -62.93962, -71.0744, 
    -68.88454, -58.6271, -43.77182, -25.82502, -8.515169, 1.41453, -2.368785, 
    -16.09882, -25.22123, -21.95242, -13.36202, -6.42433, -1.704176,
  1.099235, 0.1059141, -9.310223, -28.27311, -51.61053, -71.26639, -82.26917, 
    -80.73558, -69.13644, -51.43256, -29.62326, -7.984031, 6.05649, 4.383249, 
    -10.43218, -21.25716, -17.70652, -9.226555, -3.802008, -0.8000612,
  1.392344, 0.7480459, -9.067308, -29.56254, -55.3713, -77.64397, -90.55849, 
    -89.2873, -76.33993, -56.38977, -31.98525, -7.634667, 9.150364, 9.341149, 
    -5.745224, -17.80234, -14.59309, -6.418497, -1.957943, -0.1543795,
  1.270931, 0.3307223, -9.943935, -31.10905, -57.62258, -80.21581, -93.43466, 
    -92.22561, -78.72487, -57.98168, -32.75768, -7.616096, 9.93219, 10.65306, 
    -4.449306, -16.7849, -13.76281, -5.523272, -1.1205, 0.1760685,
  0.6025711, -1.503623, -12.41014, -33.33717, -58.60773, -79.00223, 
    -90.61551, -89.17287, -76.09286, -56.18629, -32.0011, -8.051064, 
    8.097018, 7.722486, -7.171949, -18.51095, -15.184, -6.403441, -1.203068, 
    0.2194836,
  -0.7650037, -5.226232, -17.31045, -37.58155, -60.35472, -77.08563, 
    -85.49493, -82.77731, -70.16191, -51.88966, -30.10498, -9.047067, 
    4.025129, 1.961297, -11.5921, -20.60812, -16.7964, -7.678529, -1.62451, 
    0.1317757,
  -2.893306, -11.07937, -25.26489, -45.21522, -65.5331, -79.12361, -83.99933, 
    -78.70675, -65.56998, -48.16736, -28.48831, -10.31371, 0.1995764, 
    -1.865184, -12.29841, -18.71521, -15.3679, -7.466167, -1.766869, 
    0.03671169,
  -5.563169, -18.49177, -35.63492, -56.03643, -74.95755, -87.22968, 
    -89.50784, -81.12296, -66.57057, -48.51377, -28.89139, -11.07216, 
    0.03975344, 0.9522429, -5.378934, -10.4174, -9.5241, -5.288994, 
    -1.770537, -0.1994241,
  -8.524515, -26.7611, -47.38257, -68.748, -86.85403, -98.36293, -98.97972, 
    -88.17433, -71.92631, -52.24655, -30.91523, -10.94845, 3.518342, 
    9.217065, 6.936301, 1.825674, -1.864677, -3.09588, -2.468323, -0.809729,
  -9.249249, -29.17929, -51.96335, -75.88305, -96.93556, -111.3254, 
    -117.8288, -113.9185, -98.51812, -74.46444, -45.80542, -17.94, 2.942647, 
    12.23932, 10.21183, 2.534176, -4.226498, -6.844153, -5.665792, -2.180382,
  -12.6664, -38.9888, -66.61058, -92.73451, -113.2913, -125.5022, -130.2048, 
    -124.5828, -106.6857, -79.72237, -47.80889, -16.15347, 9.230577, 
    23.25605, 24.49126, 16.43879, 4.930954, -2.612468, -3.880269, -1.75585,
  -14.57328, -44.65706, -75.54688, -103.6614, -124.5686, -135.8021, 
    -139.1838, -131.9383, -111.9728, -82.81131, -48.64419, -14.58801, 
    13.37662, 29.85775, 32.69293, 24.5848, 11.07309, 1.15343, -1.77504, 
    -1.092975,
  -15.56928, -45.46327, -71.71556, -92.39159, -106.4686, -113.7221, 
    -114.7162, -107.4785, -90.80244, -66.73724, -38.08507, -8.362162, 
    18.37354, 38.22044, 48.44943, 48.28054, 38.99044, 26.03427, 14.34644, 
    4.460615,
  -13.46367, -39.65184, -63.42309, -82.91951, -96.6851, -104, -105.5397, 
    -99.45943, -84.44608, -62.59158, -36.66788, -10.05748, 13.4709, 30.51631, 
    39.00027, 38.66381, 30.81509, 20.4518, 11.43646, 3.591021,
  -10.14759, -30.44039, -50.15623, -67.6678, -80.93779, -88.42246, -90.91759, 
    -86.76356, -74.43031, -56.07423, -34.4557, -12.79751, 5.554121, 17.97975, 
    23.4397, 22.55583, 16.81095, 10.59569, 6.080481, 1.934089,
  -6.380465, -19.85355, -34.63814, -49.56831, -62.17661, -69.98592, 
    -73.62312, -71.66872, -62.49833, -48.31501, -31.8933, -16.32005, 
    -4.450696, 2.094366, 3.647354, 2.028199, -0.9915862, -2.053634, 
    -1.028841, -0.321677,
  -2.628299, -9.167864, -18.66433, -30.6499, -42.53973, -50.99547, -55.793, 
    -55.80341, -49.79579, -39.96378, -29.14213, -20.36199, -15.96947, 
    -16.31465, -19.20486, -21.27431, -20.56582, -15.75879, -8.899869, 
    -2.851683,
  0.8756933, 0.9034257, -3.433444, -12.54638, -23.9993, -33.65077, -39.49481, 
    -40.80064, -37.48116, -31.62261, -26.28167, -24.67899, -28.70462, 
    -36.88296, -44.18758, -45.41243, -39.16687, -27.92608, -15.81563, 
    -5.050069,
  0.8911015, 1.24961, -2.114183, -9.77948, -19.82748, -29.15952, -35.2454, 
    -34.52682, -28.50697, -21.57892, -16.38186, -15.21531, -19.67405, 
    -28.48539, -36.61234, -39.14685, -35.67809, -26.41422, -14.9717, -4.693082,
  1.930065, 4.196919, 2.039731, -5.83953, -17.72589, -29.65878, -38.53556, 
    -39.71173, -33.94689, -26.07445, -18.89114, -15.72032, -20.15363, 
    -31.52027, -41.85365, -43.05293, -35.12379, -23.51552, -12.60298, 
    -3.796846,
  2.554837, 5.960961, 4.416339, -4.046748, -18.05643, -33.11748, -45.23391, 
    -48.34537, -42.56365, -33.00417, -22.49718, -15.31721, -17.2934, 
    -29.46714, -41.84047, -42.86199, -32.12576, -19.4477, -9.810641, -2.800544,
  2.969107, 7.113979, 5.877668, -3.277278, -19.31927, -37.34304, -52.62727, 
    -57.64417, -51.59405, -39.96477, -25.90501, -14.47744, -13.11626, 
    -24.88465, -39.00441, -40.82277, -29.02919, -16.08405, -7.557834, 
    -2.007024,
  3.063881, 7.354185, 6.030514, -3.778191, -21.21778, -41.01578, -58.37401, 
    -64.71446, -58.17691, -44.77964, -28.16614, -13.8526, -9.979831, 
    -20.99634, -36.13913, -38.78022, -26.86213, -13.90362, -5.981191, 
    -1.436091,
  2.754406, 6.464676, 4.644069, -5.581793, -23.30062, -42.956, -60.44616, 
    -67.11856, -60.29649, -46.27747, -28.93423, -13.91844, -9.504055, 
    -20.35887, -35.62888, -38.31065, -26.46696, -13.34204, -5.305254, 
    -1.156041,
  1.93947, 4.163197, 1.311181, -9.148438, -26.04232, -43.76116, -59.22233, 
    -64.82303, -57.87618, -44.4762, -28.33918, -14.95778, -12.18536, 
    -23.50801, -37.71339, -39.31475, -27.48147, -14.10176, -5.460116, 
    -1.160477,
  0.5221869, 0.1420009, -4.549636, -15.47872, -31.15209, -46.36754, 
    -58.43725, -61.32578, -53.67735, -41.12464, -27.18487, -16.84447, 
    -16.58522, -27.70963, -39.43091, -39.39915, -27.94717, -14.92571, 
    -5.98706, -1.341752,
  -1.448708, -5.515683, -13.01394, -25.15513, -40.22595, -53.9155, -62.69244, 
    -61.85449, -52.59767, -39.88112, -27.11827, -18.59274, -18.90531, 
    -27.74991, -36.3021, -35.49995, -25.70659, -14.57593, -6.485618, -1.625538,
  -3.621131, -11.85903, -22.82955, -37.06231, -52.70402, -66.38745, 
    -72.87751, -68.35483, -56.95993, -42.79883, -28.96911, -19.09915, 
    -16.60932, -21.24379, -26.98056, -27.07019, -20.69486, -13.23226, 
    -7.169695, -2.116976,
  -5.684139, -17.99162, -32.57747, -49.23857, -65.8384, -79.69777, -84.82082, 
    -77.68465, -64.11469, -47.8424, -31.5607, -18.36984, -11.3076, -11.14789, 
    -14.66843, -16.86762, -15.55273, -12.80096, -8.808487, -3.013565,
  -5.553138, -18.39517, -35.2719, -55.63038, -76.04054, -91.99048, -100.2877, 
    -98.3813, -86.35079, -67.73587, -47.16884, -29.72492, -19.80357, 
    -18.74048, -23.16608, -27.02344, -26.12742, -21.09965, -13.75536, 
    -4.775731,
  -7.85326, -25.38582, -46.72017, -70.18066, -91.3531, -105.828, -112.5126, 
    -108.7933, -94.05531, -72.46056, -48.64766, -27.49708, -13.47669, 
    -8.736699, -11.38696, -16.57688, -20.25335, -19.0056, -12.91293, -4.594741,
  -9.058386, -29.26061, -53.59446, -79.61563, -101.9284, -115.8013, 
    -121.1609, -115.6693, -98.70833, -74.88895, -48.93845, -25.68675, 
    -9.670026, -3.345449, -5.212833, -10.7039, -15.97189, -16.28988, 
    -11.17805, -4.005559,
  -11.65638, -34.96076, -57.55361, -77.47466, -92.31907, -100.3525, 
    -101.8497, -95.51403, -81.09953, -61.59667, -40.15944, -19.88676, 
    -3.592886, 6.841378, 11.08557, 10.16059, 5.470749, 1.066402, -0.5385838, 
    -0.4374809,
  -10.23587, -30.73641, -50.76056, -68.7275, -82.55068, -90.53269, -92.97878, 
    -88.38649, -76.10276, -58.9459, -39.96095, -22.09881, -7.903712, 
    1.100817, 4.843235, 4.341036, 0.7743988, -2.076647, -2.190695, -0.9417063,
  -7.741118, -23.4152, -39.21004, -54.10577, -66.39706, -74.33151, -78.22086, 
    -76.34232, -67.47353, -54.17206, -39.32764, -25.6558, -15.23303, 
    -8.945151, -6.350544, -6.294289, -7.847557, -7.811984, -5.190139, -1.85146,
  -4.564417, -14.12491, -24.61928, -35.69704, -46.09177, -53.96824, 
    -59.37244, -60.51036, -55.80288, -47.45165, -38.15435, -30.30528, 
    -25.28463, -23.00445, -22.19263, -21.36264, -19.84808, -15.71424, 
    -9.417927, -3.150389,
  -1.082582, -3.919825, -8.526241, -15.29177, -23.49872, -31.31873, 
    -37.88291, -41.59276, -41.25151, -38.60339, -36.16508, -35.9287, 
    -38.21638, -41.38396, -42.8317, -40.61935, -34.57825, -25.24998, 
    -14.7196, -4.814664,
  2.275205, 5.973268, 7.211608, 4.854574, -1.031033, -8.761615, -15.73113, 
    -20.91463, -24.60003, -27.92169, -33.39771, -42.66781, -54.38922, 
    -64.25104, -67.63327, -62.49702, -50.01244, -34.71252, -20.07169, 
    -6.504864,
  2.616452, 7.404431, 10.66466, 11.05412, 7.560528, -0.1264353, -9.387877, 
    -14.63397, -15.42309, -15.88454, -19.46778, -28.0617, -40.24048, 
    -51.09635, -55.60254, -52.33841, -43.21018, -31.25134, -18.54028, 
    -6.014587,
  3.556428, 10.26395, 15.40333, 17.2734, 14.52509, 6.971049, -3.910941, 
    -12.05933, -14.53053, -15.73159, -19.98103, -30.48216, -46.22049, 
    -60.21404, -64.79642, -58.45675, -45.32075, -30.89162, -17.4411, -5.5073,
  3.970726, 11.61378, 17.83783, 20.63368, 18.17886, 10.04887, -3.039524, 
    -14.23843, -18.19416, -19.15473, -21.86645, -31.09772, -47.66218, 
    -63.71815, -68.81841, -60.62263, -44.57174, -28.96491, -15.92048, 
    -4.938177,
  4.077424, 12.04651, 18.78969, 22.06576, 19.62354, 10.75359, -4.518965, 
    -18.6844, -23.97278, -24.16501, -24.23397, -30.46128, -46.05907, 
    -63.38792, -69.47752, -60.69009, -43.2392, -27.21714, -14.6776, -4.491902,
  3.848287, 11.47177, 18.10955, 21.43624, 18.98435, 9.965873, -6.47052, 
    -22.66867, -28.76331, -28.15175, -26.07715, -29.85424, -44.32526, 
    -62.27014, -69.09979, -60.22222, -42.41894, -26.25451, -13.87264, -4.19026,
  3.298074, 9.935863, 15.88343, 18.89636, 16.53082, 8.09721, -7.917347, 
    -24.25119, -30.30964, -29.41442, -26.97052, -30.50275, -44.92352, 
    -62.81638, -69.38698, -60.24179, -42.57316, -26.31895, -13.71234, -4.10881,
  2.449733, 7.495212, 12.16276, 14.41884, 12.00536, 4.294983, -10.03036, 
    -24.27971, -29.22262, -28.43768, -27.33064, -32.71125, -47.888, 
    -64.74054, -69.93749, -60.35896, -43.11366, -26.99804, -14.15318, 
    -4.261778,
  1.357289, 4.265841, 6.999104, 7.795969, 4.655156, -3.151867, -15.58109, 
    -26.25911, -29.08549, -27.98801, -28.23876, -35.30376, -50.23485, 
    -64.86404, -68.46062, -59.06521, -42.77559, -27.45614, -14.89056, 
    -4.578614,
  0.1885731, 0.6720126, 0.8683467, -0.7167377, -5.754605, -15.03493, 
    -26.28053, -33.0986, -33.21017, -30.71205, -30.42595, -36.49656, 
    -48.75221, -60.34883, -63.12164, -55.21353, -40.81245, -27.24176, 
    -15.69089, -4.995541,
  -0.7390254, -2.406255, -4.97494, -9.719902, -17.8098, -29.69583, -40.72678, 
    -44.24362, -41.35209, -36.32745, -33.35008, -35.71409, -43.40432, 
    -51.71279, -54.48349, -49.19088, -37.737, -26.78519, -16.71013, -5.560943,
  -1.309318, -4.537948, -9.576395, -17.47294, -28.72691, -43.17373, 
    -54.82326, -56.28055, -50.47813, -42.44215, -35.92974, -33.76985, 
    -36.6109, -41.82664, -44.92057, -42.78097, -35.32808, -27.5121, 
    -18.63442, -6.476995,
  -0.212682, -2.238793, -8.465997, -19.88518, -35.2553, -51.2723, -63.18666, 
    -67.96104, -65.86153, -59.89546, -54.70288, -54.09476, -58.92412, 
    -66.08591, -70.21382, -67.13058, -55.99076, -41.34515, -25.82319, 
    -8.778759,
  -1.431044, -6.119433, -15.4021, -29.80003, -47.1475, -63.40472, -75.14541, 
    -78.70289, -73.67874, -64.42246, -55.82418, -51.6784, -53.21273, 
    -58.12755, -61.80026, -60.41846, -53.26582, -41.23716, -25.91982, 
    -8.864281,
  -2.144717, -8.44824, -19.75275, -36.35234, -55.35678, -71.9381, -83.14522, 
    -85.29158, -78.00906, -66.46413, -55.85478, -50.07736, -50.44025, 
    -54.63915, -57.9654, -56.74901, -50.76525, -39.70359, -24.80021, -8.466715,
  -8.123829, -24.89276, -42.45262, -59.46831, -73.54082, -82.40317, 
    -85.87235, -82.5491, -72.27242, -58.27056, -43.71992, -31.2626, 
    -22.63214, -18.15732, -16.73889, -16.80021, -17.49954, -15.90676, 
    -10.76316, -3.838174,
  -7.21089, -22.00861, -37.36195, -52.26459, -64.88276, -73.3484, -77.63928, 
    -76.109, -68.06355, -56.38126, -44.00601, -33.37566, -26.0123, -22.12238, 
    -20.68958, -20.3441, -20.37073, -17.8855, -11.85297, -4.18349,
  -5.472926, -16.68378, -28.34984, -39.94862, -50.3663, -58.21468, -63.67735, 
    -64.88289, -60.42769, -52.62975, -44.05959, -36.81148, -32.01023, 
    -29.55377, -28.39645, -27.34754, -25.87075, -21.45788, -13.70822, 
    -4.744988,
  -3.054403, -9.402881, -16.33381, -23.87864, -31.65005, -38.73738, 
    -45.30975, -49.52071, -49.5277, -46.89065, -43.67007, -41.45502, 
    -40.71447, -40.73596, -40.20298, -37.99734, -33.83991, -26.38057, 
    -16.24769, -5.503882,
  -0.1531041, -0.7492734, -2.242223, -5.242364, -10.05993, -16.2711, 
    -23.41802, -30.10832, -34.96228, -38.60562, -42.4761, -47.43131, 
    -52.79755, -56.65681, -57.02077, -52.82568, -44.32323, -32.63549, 
    -19.61725, -6.533677,
  2.818617, 8.103104, 12.16543, 13.86491, 12.24086, 7.194193, 0.5755825, 
    -7.264355, -16.82758, -27.64317, -40.51531, -55.2969, -69.23163, 
    -78.10267, -78.88074, -71.08952, -56.25278, -39.39222, -23.38341, 
    -7.703618,
  3.198469, 9.632055, 15.76032, 20.30328, 21.25471, 16.40005, 7.298001, 
    -1.131596, -7.460329, -14.20121, -24.02783, -37.65209, -51.94029, 
    -61.65254, -63.48654, -57.75586, -46.51804, -33.85168, -20.78579, 
    -6.894806,
  4.05884, 12.29158, 20.36662, 26.92692, 29.90001, 27.14477, 18.08588, 
    6.900761, -2.061498, -11.119, -23.90399, -42.0104, -61.10789, -73.23033, 
    -73.90123, -64.81573, -50.52947, -35.35331, -20.57751, -6.646956,
  4.394483, 13.4372, 22.62601, 30.538, 34.89582, 33.37333, 23.745, 9.72751, 
    -1.543647, -11.63758, -24.82018, -44.27549, -65.95946, -79.81746, 
    -79.82101, -68.35838, -51.62528, -35.19343, -20.04989, -6.400794,
  4.384978, 13.55087, 23.18682, 31.82967, 36.99174, 36.10429, 25.74867, 
    9.172166, -4.14619, -14.53172, -26.39085, -44.76926, -67.17439, 
    -82.29577, -82.28689, -69.64839, -51.63188, -34.73534, -19.63439, 
    -6.240278,
  4.042556, 12.65691, 22.06552, 30.83534, 36.39159, 36.09589, 25.62008, 
    7.558913, -7.015485, -17.37973, -27.90048, -44.93975, -67.33202, 
    -83.10796, -83.14627, -70.01365, -51.67809, -34.63851, -19.46325, 
    -6.169725,
  3.462915, 11.02765, 19.67274, 28.05375, 33.61755, 33.74372, 23.87308, 
    6.145575, -8.316051, -18.61074, -29.12026, -46.2326, -68.58765, 
    -84.03708, -83.62164, -70.25907, -52.09925, -35.06538, -19.70615, 
    -6.252796,
  2.770844, 9.005307, 16.47991, 23.95126, 28.92234, 28.68798, 19.53753, 
    3.813135, -9.141066, -19.12549, -30.57206, -48.61253, -70.43632, 
    -84.51141, -83.37076, -70.1731, -52.42512, -35.6574, -20.32304, -6.499515,
  2.098509, 6.929605, 12.88692, 18.78885, 22.20358, 20.26703, 11.15519, 
    -1.874583, -12.45467, -21.36783, -32.87744, -50.47274, -70.30663, 
    -82.47996, -81.17667, -68.99141, -51.96763, -35.92043, -21.08793, 
    -6.847643,
  1.597559, 5.195212, 9.375569, 12.94147, 13.59787, 8.542377, -1.564678, 
    -12.10542, -19.84888, -26.49085, -35.88878, -50.44679, -66.68595, 
    -76.92629, -76.35955, -66.17456, -50.46576, -35.70988, -21.84217, 
    -7.241798,
  1.446489, 4.321128, 6.751731, 7.426328, 4.332363, -4.798001, -16.83186, 
    -25.52497, -30.10884, -33.36359, -38.85496, -48.6435, -60.48693, 
    -68.87001, -69.49727, -61.92434, -48.28355, -35.39009, -22.72446, 
    -7.725789,
  1.61335, 4.347963, 5.461213, 3.467093, -3.324752, -16.456, -31.13551, 
    -39.0507, -40.5266, -40.01397, -41.16863, -46.05663, -53.67211, 
    -60.29277, -62.08591, -57.36759, -46.68387, -36.1116, -24.40054, -8.519246,
  3.023952, 7.744618, 8.741632, 4.356828, -5.72777, -19.9312, -33.78089, 
    -44.40368, -51.652, -56.86316, -63.40041, -73.3382, -85.18733, -94.4179, 
    -96.37325, -88.80106, -72.29034, -52.81692, -32.92555, -11.18976,
  2.20064, 5.151244, 4.10149, -2.517782, -14.63045, -30.03822, -45.1216, 
    -55.53382, -60.00438, -61.69787, -64.6406, -71.1255, -80.11458, 
    -87.66558, -89.51073, -83.62299, -70.8148, -53.53746, -33.48895, -11.42641,
  1.606989, 3.323234, 0.9024963, -7.236497, -20.7752, -36.94976, -52.32231, 
    -61.98739, -64.43795, -63.89883, -64.94531, -70.06125, -78.17312, 
    -85.13405, -86.57526, -80.77093, -69.09129, -52.65952, -32.81218, 
    -11.18748,
  -4.393363, -13.91285, -25.04863, -37.38087, -49.32267, -58.7972, -65.24299, 
    -66.75474, -62.67393, -55.96154, -49.46942, -45.13558, -43.50741, 
    -43.60228, -43.5568, -41.94547, -38.69165, -31.69678, -20.45307, -7.103701,
  -3.841769, -12.08922, -21.58786, -32.07109, -42.4381, -51.15933, -58.02564, 
    -61.04413, -59.04088, -54.46587, -49.78609, -46.68896, -45.63744, 
    -45.79066, -45.57798, -43.76413, -40.21685, -32.77583, -21.0613, -7.298522,
  -2.740978, -8.582199, -15.2599, -22.76578, -30.6698, -38.1785, -45.55211, 
    -50.8325, -52.20479, -51.28609, -49.90757, -49.32095, -49.76505, 
    -50.46976, -50.16209, -47.82681, -43.30015, -34.67952, -22.01452, 
    -7.577494,
  -1.106576, -3.50845, -6.442348, -10.22697, -15.13424, -21.14174, -28.79078, 
    -36.49289, -42.14302, -46.23557, -49.70756, -53.14069, -56.30362, 
    -58.27517, -57.94158, -54.49452, -47.85049, -37.15695, -23.18885, 
    -7.901182,
  1.035652, 3.014304, 4.571929, 5.028873, 3.464279, -0.8352041, -8.103207, 
    -17.6455, -28.10709, -38.62361, -48.94469, -58.59924, -66.36488, 
    -70.67065, -70.30029, -64.73299, -54.25732, -40.40097, -24.82189, -8.36698,
  3.400896, 10.15442, 16.49191, 21.42615, 23.51356, 21.37622, 15.80647, 
    5.8869, -9.491047, -27.99202, -47.8065, -66.72659, -81.48663, -89.03216, 
    -87.96559, -78.63055, -62.30893, -44.27247, -26.90214, -8.984812,
  3.619931, 11.17078, 19.16957, 26.56473, 31.04361, 29.33701, 21.87587, 
    11.66472, -0.02813339, -13.54054, -29.43339, -46.58674, -61.1315, 
    -69.00449, -68.78599, -61.6268, -49.15998, -36.1959, -22.88437, -7.724791,
  4.342945, 13.43081, 23.21555, 32.79996, 40.12821, 42.18237, 36.69694, 
    24.65352, 9.69413, -8.030391, -29.37633, -52.87489, -72.32845, -81.53502, 
    -79.38799, -69.14564, -54.81794, -39.34536, -23.43853, -7.688281,
  4.634141, 14.42992, 25.24652, 36.30029, 45.65899, 50.46533, 46.33804, 
    32.55487, 14.96348, -5.427986, -29.83402, -57.33242, -80.23746, 
    -90.35184, -86.63659, -73.92656, -57.88743, -41.0067, -23.85275, -7.733884,
  4.598764, 14.44386, 25.61343, 37.40118, 47.90788, 54.3117, 51.00439, 
    35.94065, 16.30775, -5.589627, -30.86843, -59.78784, -84.47476, 
    -95.18694, -90.55932, -76.39411, -59.30996, -41.85257, -24.23952, 
    -7.844551,
  4.267803, 13.55441, 24.43075, 36.26593, 47.1888, 54.40755, 51.79908, 
    36.37379, 15.70065, -6.913568, -32.22311, -61.33544, -86.63574, 
    -97.50867, -92.33871, -77.51321, -60.1125, -42.4887, -24.64871, -7.988968,
  3.805552, 12.23106, 22.41286, 33.77518, 44.44677, 51.56135, 49.33023, 
    34.6019, 14.21407, -8.442529, -33.93956, -63.08534, -88.07612, -98.46351, 
    -92.93845, -78.03021, -60.65265, -43.07847, -25.19561, -8.204498,
  3.409904, 11.02827, 20.3676, 30.84521, 40.51883, 46.25386, 43.49106, 
    29.941, 10.82434, -11.09658, -36.3783, -64.76332, -88.32384, -97.83748, 
    -92.46395, -78.0949, -60.78038, -43.4561, -25.86182, -8.494976,
  3.227986, 10.34169, 18.81831, 27.96648, 35.71624, 38.61873, 34.0194, 
    21.35798, 4.003095, -16.10452, -39.50568, -65.22916, -86.21291, 
    -94.95685, -90.5693, -77.44975, -60.29007, -43.461, -26.51818, -8.81583,
  3.329624, 10.35568, 17.99166, 25.30851, 30.11415, 28.89013, 21.21936, 
    8.846887, -6.298627, -23.25243, -42.75172, -63.9972, -81.62752, 
    -89.76849, -86.9576, -75.67271, -59.08052, -43.10473, -27.08496, -9.134712,
  3.752707, 11.20684, 18.16818, 23.33654, 24.44465, 18.2999, 6.662737, 
    -6.000495, -18.43988, -31.17101, -45.56675, -61.56718, -75.59433, 
    -83.06039, -81.84438, -72.65413, -57.28385, -42.63876, -27.6944, -9.50054,
  4.394787, 12.72132, 19.43776, 22.79116, 20.36811, 9.372334, -6.819064, 
    -20.53815, -30.16805, -38.40879, -47.67952, -58.71175, -69.33855, 
    -75.97927, -76.10863, -69.15381, -55.84414, -42.99904, -28.96526, 
    -10.13062,
  5.936816, 16.72962, 24.31616, 26.69468, 22.38387, 11.20421, -3.489571, 
    -19.83211, -37.51689, -55.31067, -73.85651, -92.75522, -108.8971, 
    -117.981, -117.0803, -105.651, -85.02433, -61.93663, -38.65374, -13.14887,
  5.37873, 15.02945, 21.38612, 22.35267, 16.38197, 3.48975, -13.72486, 
    -31.17101, -46.56936, -60.71054, -75.42812, -90.86839, -104.3943, 
    -112.0836, -111.2243, -101.4642, -84.34222, -63.18384, -39.54494, 
    -13.49674,
  4.870243, 13.55093, 19.02599, 19.12522, 12.20812, -1.549017, -19.76282, 
    -37.32125, -51.20947, -63.34369, -76.31356, -90.50851, -103.1616, 
    -110.135, -108.7731, -99.12516, -83.18954, -62.83075, -39.2463, -13.3956,
  1.033209, 2.333178, 1.551694, -2.130917, -8.902002, -18.08384, -29.34687, 
    -40.04281, -47.98064, -54.55259, -61.09607, -67.93031, -74.07926, 
    -77.77001, -77.4638, -72.73531, -64.39781, -50.97495, -32.44783, -11.18091,
  1.279617, 3.14831, 3.142706, 0.4903879, -5.123552, -13.36937, -24.33741, 
    -35.65025, -44.90605, -52.93937, -60.58683, -67.94698, -74.16681, 
    -77.79751, -77.54313, -72.95021, -64.62053, -51.08442, -32.47045, 
    -11.17731,
  1.74343, 4.686269, 6.12693, 5.32695, 1.720301, -4.921885, -15.25489, 
    -27.45085, -38.95488, -49.6689, -59.57642, -68.33776, -75.1563, 
    -78.95393, -78.75602, -74.1001, -65.32224, -51.27916, -32.45022, -11.13845,
  2.427466, 6.931817, 10.40231, 12.09958, 11.12362, 6.571548, -2.634064, 
    -15.60443, -30.0961, -44.73613, -58.26279, -69.58961, -77.7823, 
    -82.04905, -81.74166, -76.4531, -66.32269, -51.24947, -32.22029, -11.01061,
  3.430719, 10.13881, 16.27049, 21.04565, 23.20536, 21.14231, 13.83768, 
    0.7135119, -17.40026, -37.59321, -56.81753, -72.67333, -83.62393, 
    -88.88723, -88.10271, -81.10722, -68.08984, -51.20005, -31.98344, 
    -10.87303,
  4.683819, 14.07267, 23.29539, 31.56645, 37.37519, 38.51014, 34.53864, 
    22.67613, 0.4845467, -27.62013, -55.85261, -79.28648, -94.86622, 
    -101.4858, -99.30315, -88.95977, -71.15765, -51.51197, -31.99999, 
    -10.81817,
  4.31409, 13.3056, 22.98009, 32.61176, 40.16185, 42.16043, 38.00666, 
    27.4301, 9.756756, -12.69861, -36.11147, -56.38877, -70.159, -75.96087, 
    -74.24423, -66.29124, -52.95126, -39.68956, -25.79582, -8.847259,
  4.633805, 14.39563, 25.25812, 36.89625, 47.87291, 55.24245, 55.51594, 
    45.20393, 24.28806, -4.838494, -36.63816, -64.20035, -81.74329, 
    -87.51693, -83.62975, -73.61917, -60.16718, -44.55865, -27.19328, 
    -9.045411,
  4.819368, 15.04645, 26.66807, 39.64137, 53.0362, 64.62175, 68.66144, 
    58.9219, 35.98495, 1.72841, -37.27608, -71.39281, -92.15408, -97.58286, 
    -91.55965, -79.59859, -65.83797, -48.55535, -28.68588, -9.399423,
  4.857599, 15.21107, 27.11109, 40.66113, 55.22345, 69.04173, 75.498, 
    66.75526, 43.03105, 5.638513, -38.2446, -76.85983, -99.5955, -104.4773, 
    -96.8475, -83.49248, -69.13383, -50.98096, -29.93661, -9.785913,
  4.755974, 14.91742, 26.66111, 40.13842, 54.81551, 69.06302, 76.51183, 
    68.85981, 45.17179, 6.436099, -39.7313, -80.32958, -103.7194, -108.109, 
    -99.63966, -85.59659, -70.62227, -52.15308, -30.83906, -10.1185,
  4.699801, 14.70823, 26.18702, 39.23683, 53.24988, 66.37254, 73.27747, 
    66.19881, 42.73426, 4.00596, -41.98885, -82.09612, -105.0266, -109.2551, 
    -100.8268, -86.68864, -70.96487, -52.45655, -31.46747, -10.39799,
  4.883609, 15.14827, 26.57396, 39.09414, 51.86219, 62.55, 67.27346, 59.5859, 
    36.00756, -1.613823, -45.0867, -82.45098, -104.077, -108.6346, -101.1204, 
    -87.34691, -70.68727, -52.2399, -31.92446, -10.64338,
  5.373857, 16.4269, 28.10243, 40.03043, 50.98701, 58.11239, 59.07687, 
    49.40555, 25.55061, -9.69908, -48.62289, -81.62768, -101.3849, -106.5733, 
    -100.5476, -87.50648, -70.00298, -51.7305, -32.25006, -10.85628,
  6.105356, 18.35563, 30.47246, 41.64293, 50.17163, 52.80605, 48.76751, 
    36.17043, 12.51938, -18.99515, -52.07589, -79.96073, -97.46117, 
    -103.1192, -98.63361, -86.58204, -68.74162, -50.95934, -32.43462, 
    -11.03349,
  7.007501, 20.74608, 33.43989, 43.72357, 49.38328, 46.98205, 37.17217, 
    21.21628, -1.444974, -28.2628, -55.10248, -77.81262, -92.80983, 
    -98.46067, -95.17116, -84.23648, -66.79745, -49.99356, -32.55529, 
    -11.21131,
  7.999888, 23.43508, 36.96716, 46.62938, 49.58723, 42.17392, 26.20689, 
    6.580547, -14.65386, -36.50075, -57.38296, -75.29906, -87.78883, 
    -93.09442, -90.74448, -81.13076, -64.87763, -49.49514, -33.09093, 
    -11.56331,
  9.577853, 27.82061, 43.26578, 53.80897, 57.15192, 51.26511, 37.37611, 
    14.69838, -17.49131, -53.70173, -88.42303, -116.9376, -135.5744, 
    -142.437, -137.4842, -121.8274, -97.11593, -70.57229, -44.05771, -14.99034,
  9.307986, 27.04134, 42.02894, 52.0355, 54.4099, 46.77795, 29.3104, 
    3.735563, -27.37374, -60.0256, -90.55293, -115.4218, -131.5346, 
    -137.1944, -132.4471, -118.4894, -97.00711, -72.10725, -45.13902, 
    -15.40201,
  8.944462, 26.03051, 40.56985, 50.31192, 52.40186, 44.22452, 25.32287, 
    -1.495798, -32.20142, -63.51608, -92.52141, -116.0101, -130.9068, 
    -135.5742, -130.309, -116.6232, -96.40084, -72.23292, -45.18472, -15.42421,
  4.291628, 12.08061, 17.57837, 19.43825, 16.53013, 8.405453, -5.322376, 
    -22.01695, -38.42069, -54.22458, -69.03322, -81.84467, -91.14249, 
    -95.49011, -94.17179, -87.46886, -76.48921, -59.96138, -38.02742, 
    -13.07415,
  4.408135, 12.45476, 18.29593, 20.66093, 18.45312, 11.1004, -2.03755, 
    -18.68699, -35.64581, -52.21315, -67.5972, -80.66148, -90.04453, 
    -94.54194, -93.51149, -87.09694, -76.20406, -59.66778, -37.79865, 
    -12.98442,
  4.599088, 13.11471, 19.67056, 23.10155, 22.28907, 16.37756, 4.369128, 
    -12.15151, -30.22874, -48.45076, -65.29601, -79.28668, -89.16901, 
    -94.02921, -93.35852, -87.14165, -75.99065, -59.18914, -37.38988, 
    -12.81773,
  4.841351, 13.9945, 21.592, 26.58448, 27.76622, 23.85856, 13.609, -2.478992, 
    -22.19806, -43.10767, -62.55251, -78.40014, -89.34563, -94.74123, 
    -94.25772, -87.77631, -75.6299, -58.21584, -36.63741, -12.5224,
  5.239607, 15.38754, 24.4871, 31.59839, 35.37868, 34.0261, 26.36916, 
    11.33438, -10.63862, -35.82824, -59.83157, -79.24934, -92.32377, 
    -98.52416, -97.76431, -90.02676, -75.54971, -56.92306, -35.70738, -12.163,
  5.801224, 17.29268, 28.30613, 38.05888, 45.14075, 47.26981, 43.63743, 
    30.88551, 6.023689, -26.04205, -58.01484, -83.85239, -100.5589, 
    -107.6293, -105.5775, -95.02443, -76.4939, -55.81719, -34.90278, -11.84142,
  4.929628, 15.01929, 25.50104, 35.74799, 44.05672, 47.3457, 44.77966, 
    34.59041, 14.83735, -11.38081, -38.05648, -59.69138, -73.42171, 
    -78.92855, -77.15992, -69.22746, -55.69695, -42.13008, -27.57698, 
    -9.501319,
  4.865362, 15.00805, 26.11567, 38.07051, 49.8611, 58.96608, 61.76062, 
    53.01761, 30.59848, -2.771219, -38.41836, -67.02171, -83.73692, 
    -88.83274, -85.22191, -76.07301, -63.32386, -47.61897, -29.38644, 
    -9.832579,
  4.906175, 15.22386, 26.81608, 39.91149, 54.12665, 67.82905, 75.22348, 
    68.14595, 44.35244, 5.113962, -39.03772, -74.48814, -93.86401, -98.19686, 
    -92.60117, -82.1629, -70.06203, -52.6005, -31.28613, -10.29051,
  5.004813, 15.53109, 27.39042, 40.95985, 56.22287, 72.18216, 82.35201, 
    77.07654, 53.22396, 10.37782, -40.01207, -80.56976, -101.6269, -105.1122, 
    -97.97665, -86.44781, -74.09808, -55.58002, -32.74511, -10.72797,
  5.127217, 15.85175, 27.79021, 41.31536, 56.50985, 72.52337, 83.43197, 
    79.515, 56.10031, 11.81386, -41.51339, -84.4352, -106.1248, -109.1264, 
    -101.252, -88.99489, -75.66225, -56.67424, -33.6362, -11.06085,
  5.402533, 16.58007, 28.69798, 41.99442, 56.41696, 70.82943, 80.60003, 
    76.91727, 53.48021, 9.171733, -43.86568, -86.34499, -107.8636, -111.0054, 
    -103.2276, -90.52679, -75.67989, -56.51707, -34.07584, -11.29018,
  5.953161, 18.08626, 30.73994, 43.89353, 57.16275, 68.86768, 75.84261, 
    70.71365, 46.30305, 2.891491, -47.21902, -86.95144, -107.6659, -111.4804, 
    -104.482, -91.59601, -75.05613, -55.81301, -34.27365, -11.45656,
  6.769872, 20.34726, 33.88934, 46.99315, 58.77941, 66.94756, 69.67149, 
    61.42998, 35.52511, -5.927512, -51.2167, -86.73521, -106.0893, -110.6846, 
    -104.7986, -92.02396, -74.10044, -54.92442, -34.34314, -11.58364,
  7.736982, 23.0214, 37.59354, 50.55965, 60.43706, 64.383, 61.76157, 
    49.39036, 22.36061, -15.89979, -55.31268, -85.97079, -103.4391, 
    -108.4199, -103.5417, -91.15765, -72.55282, -53.81108, -34.26258, 
    -11.66703,
  8.774526, 25.8767, 41.4961, 54.17706, 61.79189, 61.09663, 52.49832, 
    35.62997, 8.296672, -25.79894, -59.01564, -84.72382, -99.9044, -104.6854, 
    -100.4794, -88.70145, -70.24565, -52.43353, -34.04543, -11.7201,
  9.849055, 28.85858, 45.64613, 58.16624, 63.5766, 58.19268, 43.35963, 
    21.90655, -5.131475, -34.59056, -61.75634, -82.78426, -95.62717, 
    -99.94283, -96.28411, -85.38674, -67.78671, -51.28521, -34.05777, 
    -11.87605,
  11.40514, 33.29311, 52.38371, 66.60625, 73.54836, 70.5857, 57.90094, 
    33.08203, -5.824669, -51.34517, -94.03875, -126.6398, -145.7503, 
    -151.1895, -144.3479, -126.9591, -100.7292, -73.01875, -45.52278, 
    -15.47534,
  11.2758, 32.92701, 51.82057, 65.7746, 72.02348, 67.4866, 51.14913, 
    22.80149, -15.80416, -58.01268, -96.36099, -125.1733, -141.769, 
    -146.1151, -139.5995, -123.9211, -100.6932, -74.46478, -46.54748, 
    -15.86514,
  11.01151, 32.19596, 50.79148, 64.64063, 70.83296, 66.00722, 48.32109, 
    18.35252, -20.52596, -61.9235, -98.88228, -126.1317, -141.2726, 
    -144.5343, -137.5681, -122.2578, -100.2712, -74.71067, -46.67527, 
    -15.91486,
  8.240132, 23.78895, 36.60862, 44.92328, 46.85691, 40.78094, 25.12977, 
    1.800361, -25.0286, -52.43294, -77.08913, -96.16417, -108.0081, 
    -112.2403, -109.3797, -100.4408, -86.7221, -67.27385, -42.45175, -14.55123,
  8.200761, 23.67164, 36.42483, 44.72748, 46.79196, 41.07082, 26.07843, 
    3.505397, -22.75589, -49.79891, -74.30717, -93.47694, -105.6729, 
    -110.449, -108.1675, -99.65762, -86.08888, -66.72372, -42.08156, -14.41693,
  8.113749, 23.45371, 36.20388, 44.72594, 47.33693, 42.50433, 28.82406, 
    7.477217, -18.249, -45.2902, -70.13487, -89.86832, -102.8151, -108.4578, 
    -106.9786, -98.94022, -85.27588, -65.84084, -41.46987, -14.1895,
  7.932757, 23.01161, 35.78388, 44.76161, 48.36425, 44.96878, 33.32206, 
    13.73478, -11.60756, -39.25453, -65.18804, -86.14045, -100.2735, 
    -106.9729, -106.2507, -98.40537, -84.09576, -64.37649, -40.48552, 
    -13.82753,
  7.734846, 22.58159, 35.57209, 45.42195, 50.63586, 49.36599, 40.61791, 
    23.38511, -2.028719, -31.5813, -60.19977, -83.72459, -99.83447, 
    -107.7408, -107.3784, -98.95007, -82.96076, -62.51997, -39.27045, 
    -13.38282,
  7.551493, 22.26143, 35.75163, 47.03446, 54.75391, 56.79501, 52.2749, 
    38.2257, 12.0057, -21.85598, -56.22065, -84.78181, -104.0561, -113.0862, 
    -112.1304, -101.7865, -82.73576, -60.84539, -38.11433, -12.94634,
  6.039618, 18.0466, 29.68441, 40.24487, 48.40165, 51.8882, 49.88479, 
    39.82293, 19.4492, -8.143042, -36.46702, -59.59697, -74.65697, -81.39113, 
    -80.62015, -73.25707, -59.90039, -45.71012, -29.85962, -10.29398,
  5.400998, 16.38728, 27.78312, 39.45786, 50.72522, 59.71841, 63.15917, 
    55.27786, 33.47567, 0.4312648, -35.08621, -63.88568, -81.4904, -88.2475, 
    -86.68092, -79.28532, -67.38486, -51.4127, -32.08335, -10.80075,
  5.134694, 15.71242, 27.09318, 39.51936, 52.89622, 66.13559, 73.99136, 
    67.89632, 45.23943, 7.62835, -34.49327, -68.57307, -88.25134, -94.56503, 
    -91.92601, -84.43081, -74.25148, -56.67662, -34.08121, -11.27323,
  5.238698, 16.02108, 27.62032, 40.39758, 54.5941, 69.7392, 79.92184, 
    75.13611, 52.23901, 11.81313, -34.76432, -72.44777, -93.41947, -99.31619, 
    -95.8709, -88.01691, -78.2238, -59.56137, -35.2856, -11.59525,
  5.630913, 17.11274, 29.17776, 42.11368, 56.21839, 71.17766, 81.63423, 
    77.64085, 54.7581, 12.97701, -35.90012, -75.53784, -97.35394, -103.2224, 
    -99.30579, -90.61707, -79.47243, -60.16187, -35.77577, -11.77814,
  6.307398, 19.011, 31.91858, 45.10567, 58.68353, 72.06361, 81.17254, 
    77.14874, 53.92542, 11.43765, -38.30432, -78.68052, -101.0027, -107.0678, 
    -102.7644, -92.74728, -79.0678, -59.34043, -35.78895, -11.86068,
  7.247163, 21.67542, 35.84733, 49.52058, 62.41668, 73.40338, 79.80676, 
    74.25948, 49.66692, 6.725833, -42.37789, -81.89275, -103.9653, -110.2057, 
    -105.6654, -94.32887, -78.00198, -58.01888, -35.59317, -11.89432,
  8.346726, 24.80242, 40.48219, 54.74113, 66.7593, 74.76543, 77.27155, 
    68.56991, 41.77993, -0.9997317, -47.71867, -84.62111, -105.4518, 
    -111.6144, -107.0242, -94.81821, -76.54202, -56.58528, -35.29667, 
    -11.89726,
  9.463017, 27.95759, 45.08916, 59.74955, 70.50594, 75.01166, 72.75079, 
    59.88408, 30.95791, -10.55888, -53.41743, -86.45353, -105.1642, 
    -110.7763, -106.1535, -93.61445, -74.39172, -54.91164, -34.81499, 
    -11.84039,
  10.53483, 30.95242, 49.3449, 64.10587, 73.19199, 73.82573, 66.33749, 
    48.98026, 18.57892, -20.49683, -58.5366, -87.09283, -103.1623, -107.8025, 
    -103.0763, -90.64445, -71.41641, -52.88129, -34.08475, -11.70427,
  11.58956, 33.89054, 53.48301, 68.23518, 75.47165, 72.04095, 59.22709, 
    37.53116, 6.327109, -29.43149, -62.20078, -86.26521, -99.75977, 
    -103.4506, -98.73998, -86.75446, -68.07923, -50.76007, -33.3191, -11.56719,
  13.06696, 38.18725, 60.29855, 77.3452, 86.96268, 86.28497, 74.98669, 
    49.8107, 7.558745, -43.75622, -92.2069, -128.3356, -148.4685, -153.4111, 
    -145.5685, -127.2639, -100.4139, -72.46733, -45.03008, -15.27581,
  13.06275, 38.15941, 60.19547, 77.0114, 85.9816, 83.91941, 69.45884, 
    40.86005, -1.683559, -50.17993, -94.39688, -126.7138, -144.4034, 
    -148.431, -141.0686, -124.4195, -100.1559, -73.48029, -45.77666, -15.56626,
  12.91217, 37.73316, 59.5735, 76.30864, 85.26282, 83.08433, 67.58598, 
    37.39128, -5.88354, -54.09324, -97.12593, -127.7841, -143.9006, 
    -146.8691, -139.1731, -122.9494, -99.80146, -73.68826, -45.87539, 
    -15.60319,
  10.04381, 29.08354, 45.06968, 56.06687, 60.03114, 55.02169, 39.07564, 
    13.59136, -17.15758, -49.17002, -77.76648, -99.29693, -112.1241, 
    -116.3526, -112.9796, -103.2802, -88.63619, -68.38164, -43.01706, 
    -14.71782,
  9.927561, 28.73908, 44.50966, 55.32632, 59.21372, 54.34459, 38.97417, 
    14.44943, -15.25373, -46.3559, -74.45477, -96.03316, -109.3632, 
    -114.3192, -111.651, -102.4465, -87.98959, -67.85217, -42.68184, -14.59955,
  9.726068, 28.17239, 43.68352, 54.41659, 58.49773, 54.18742, 40.02007, 
    17.04025, -11.4142, -41.68882, -69.55646, -91.55912, -105.819, -111.9154, 
    -110.2646, -101.6596, -87.18294, -67.03307, -42.14672, -14.40474,
  9.392424, 27.25578, 42.41954, 53.17255, 57.76731, 54.48534, 42.21141, 
    21.37917, -5.765582, -35.54113, -63.68719, -86.64382, -102.2741, -109.79, 
    -109.2271, -101.0504, -86.09441, -65.74258, -41.31156, -14.1005,
  8.989412, 26.18794, 41.08024, 52.15543, 57.80342, 56.21687, 46.63631, 
    28.49981, 2.375637, -27.8868, -57.58828, -82.65295, -100.3984, -109.5534, 
    -109.8137, -101.4505, -85.16856, -64.21549, -40.31529, -13.73328,
  8.541668, 25.0585, 39.87038, 51.77676, 59.36332, 60.6733, 54.93389, 
    40.03249, 14.27275, -18.42779, -52.22705, -81.56948, -102.583, -113.4078, 
    -113.7108, -104.022, -85.27964, -63.02293, -39.40255, -13.37391,
  6.787729, 20.08327, 32.44728, 42.99218, 50.49689, 53.24459, 50.52015, 
    39.9796, 20.31677, -5.723125, -32.96238, -56.41773, -72.91336, -81.29758, 
    -81.78583, -75.16957, -62.25743, -47.66648, -30.94455, -10.64694,
  5.884603, 17.65283, 29.3147, 40.52448, 50.57084, 57.96088, 59.88689, 
    51.34303, 31.14891, 1.966418, -29.87685, -57.61777, -76.73164, -85.98579, 
    -86.63435, -80.61966, -69.15738, -53.01039, -33.22999, -11.21943,
  5.414874, 16.3903, 27.69883, 39.32965, 51.02206, 61.82369, 67.18475, 
    59.72861, 38.92463, 7.31171, -28.03046, -58.99326, -79.86134, -89.36469, 
    -89.86311, -84.50862, -75.09183, -57.63435, -34.95753, -11.61599,
  5.43995, 16.47864, 27.89581, 39.76823, 52.07461, 64.32802, 71.22463, 
    64.05476, 42.61678, 9.572456, -27.58141, -60.18132, -81.93771, -91.54511, 
    -91.92548, -86.79817, -78.24675, -59.92287, -35.73077, -11.78173,
  5.886308, 17.74454, 29.77297, 41.96433, 54.32481, 66.51073, 73.49023, 
    66.42196, 44.44191, 10.24898, -28.3278, -62.25633, -84.88861, -94.76104, 
    -94.84996, -88.93898, -79.17713, -60.20327, -35.88361, -11.82982,
  6.688513, 20.03171, 33.19866, 45.98497, 58.23475, 69.39938, 75.46319, 
    68.3905, 45.76689, 10.01535, -30.63214, -66.37185, -90.00988, -99.95021, 
    -99.15967, -91.37981, -78.78129, -59.2374, -35.68983, -11.82405,
  7.748354, 23.06846, 37.79169, 51.42953, 63.4854, 72.94358, 77.04393, 
    69.01968, 45.01035, 7.402452, -35.03903, -71.82939, -95.65688, -105.141, 
    -103.1879, -93.3269, -77.65997, -57.74113, -35.32479, -11.79082,
  8.913647, 26.40222, 42.81145, 57.29662, 68.88569, 75.99532, 77.02196, 
    66.64888, 40.50884, 1.521152, -41.11491, -77.01403, -99.63958, -108.1535, 
    -105.2015, -93.83587, -75.9297, -56.01898, -34.82257, -11.72077,
  10.02947, 29.56151, 47.45622, 62.46127, 73.08005, 77.24005, 74.34425, 
    60.65836, 32.37604, -6.795722, -47.67559, -80.827, -101.0742, -108.2025, 
    -104.4846, -92.3685, -73.36919, -53.96436, -34.07167, -11.56863,
  11.04396, 32.38654, 51.45041, 66.54333, 75.66586, 76.43605, 69.18934, 
    51.87383, 22.02031, -15.94964, -53.50937, -82.78377, -100.0597, 
    -105.6013, -101.3025, -89.04276, -69.9539, -51.49781, -33.00114, -11.30611,
  12.01039, 35.05259, 55.12458, 70.05489, 77.34271, 74.44582, 62.83817, 
    42.16443, 11.394, -24.33, -57.68697, -82.78879, -97.21466, -101.3951, 
    -96.78726, -84.75364, -66.05378, -48.76075, -31.74498, -10.9837,
  13.40228, 39.12719, 61.66957, 78.93784, 88.6171, 87.94131, 76.95142, 
    53.08418, 13.15399, -35.96131, -83.60303, -120.4215, -141.8523, 
    -147.9215, -140.8511, -123.1658, -97.025, -69.86487, -43.32434, -14.67661,
  13.42191, 39.14464, 61.56162, 78.46664, 87.36015, 85.36028, 71.75484, 
    45.07284, 4.887927, -41.74662, -85.49105, -118.6687, -137.7457, 
    -142.9885, -136.4463, -120.3231, -96.45749, -70.45198, -43.80247, 
    -14.87345,
  13.31299, 38.8238, 61.05409, 77.8176, 86.60003, 84.45993, 70.00558, 
    41.98917, 1.172837, -45.23087, -87.92951, -119.5813, -137.1899, 
    -141.4628, -134.6439, -118.9281, -96.05155, -70.54243, -43.82304, 
    -14.88205,
  11.07763, 32.08445, 49.76069, 62.06691, 66.94547, 62.47637, 46.77023, 
    21.0636, -10.53401, -43.822, -73.78439, -96.46599, -110.0881, -114.7671, 
    -111.579, -101.8824, -87.12671, -66.9608, -42.02507, -14.35796,
  10.91444, 31.60583, 48.99416, 61.05723, 65.78718, 61.36536, 46.15677, 
    21.42759, -8.970047, -41.11256, -70.3867, -93.05024, -107.2133, 
    -112.6953, -110.2802, -101.1291, -86.59502, -66.55972, -41.79337, 
    -14.27914,
  10.65533, 30.86796, 47.88385, 59.73763, 64.50231, 60.44899, 46.28834, 
    23.1227, -5.7682, -36.68275, -65.38416, -88.33476, -103.4838, -110.2474, 
    -108.9828, -100.5271, -86.03668, -66.002, -41.45656, -14.15796,
  10.25884, 29.75541, 46.26622, 57.93574, 62.94931, 59.62976, 47.10867, 
    26.09155, -1.089865, -30.87551, -59.30752, -82.97869, -99.58135, 
    -108.0043, -108.0716, -100.2342, -85.40829, -65.18016, -40.94619, 
    -13.96982,
  9.78154, 28.44676, 44.46714, 56.15877, 61.84069, 59.8153, 49.58212, 
    31.16848, 5.58511, -23.69872, -52.78618, -78.14509, -96.95475, -107.3854, 
    -108.6848, -101.0156, -85.19452, -64.37833, -40.39397, -13.75351,
  9.241111, 27.01515, 42.67531, 54.81076, 61.92664, 62.25337, 55.16405, 
    39.60865, 15.14099, -14.98399, -46.59524, -75.45145, -97.64326, 
    -110.3366, -112.3353, -103.91, -86.2094, -64.10777, -39.96418, -13.5474,
  7.417354, 21.78325, 34.68494, 45.00953, 51.56314, 53.1651, 49.21587, 
    37.92844, 19.50529, -3.688805, -28.34317, -51.12852, -68.8548, -79.1893, 
    -81.34889, -75.84415, -63.68135, -48.85249, -31.47618, -10.80113,
  6.394558, 18.9831, 30.87771, 41.40342, 49.69753, 54.63608, 54.05248, 
    44.31673, 26.27876, 2.460468, -23.866, -49.1901, -69.48972, -81.64188, 
    -84.95628, -80.52855, -69.54009, -53.39215, -33.57085, -11.36137,
  5.771854, 17.26763, 28.50061, 39.04631, 48.30476, 55.44102, 56.93515, 
    47.56144, 29.46113, 5.572533, -21.07595, -47.30937, -68.7743, -81.82281, 
    -85.9212, -82.78267, -73.87194, -56.8233, -34.78866, -11.6191,
  5.664783, 16.982, 28.12676, 38.72336, 48.28508, 56.25462, 58.35191, 
    48.41285, 29.76459, 6.00735, -20.07848, -46.0022, -67.62964, -81.06685, 
    -85.67088, -83.34715, -75.77163, -58.24456, -35.04455, -11.6111,
  6.044202, 18.07952, 29.82053, 40.8289, 50.62264, 58.75038, 60.83088, 
    50.38479, 30.87566, 6.324297, -20.3766, -46.92781, -69.19897, -83.0211, 
    -87.53707, -84.69402, -76.4071, -58.35453, -34.94675, -11.55207,
  6.836281, 20.36931, 33.36337, 45.25328, 55.46434, 63.4212, 65.28479, 
    54.79535, 34.17796, 7.322654, -22.24612, -51.34532, -75.08795, -88.98288, 
    -92.31857, -87.36305, -76.37223, -57.62898, -34.72528, -11.50909,
  7.901481, 23.44678, 38.1188, 51.15623, 61.75698, 68.99491, 69.97796, 
    59.12569, 36.89463, 6.890922, -26.38266, -58.25244, -82.92482, -96.037, 
    -97.45007, -89.81004, -75.55573, -56.28537, -34.34401, -11.45187,
  9.047827, 26.73646, 43.12457, 57.17757, 67.74217, 73.44008, 72.45848, 
    60.24946, 35.98511, 3.263208, -32.47186, -65.32961, -89.28779, -100.7775, 
    -100.2924, -90.52452, -73.76159, -54.43027, -33.70955, -11.32861,
  10.10128, 29.7124, 47.49384, 62.07559, 71.90709, 75.24699, 71.36806, 
    56.98361, 30.83767, -3.228763, -39.2209, -70.79163, -92.5004, -101.9049, 
    -99.92021, -88.94788, -70.88253, -52.03928, -32.70998, -11.08585,
  11.0088, 32.21596, 50.96568, 65.51045, 73.93085, 74.34107, 67.10572, 
    50.27196, 22.83715, -11.01007, -45.25815, -73.90815, -92.57258, 
    -99.83725, -96.78374, -85.38347, -67.0807, -49.15706, -31.31416, -10.70161,
  11.83839, 34.46323, 53.92799, 68.05599, 74.58497, 71.73401, 61.21634, 
    42.30428, 14.207, -18.35642, -49.69819, -74.78139, -90.42021, -95.88902, 
    -92.17273, -80.76141, -62.66035, -45.84082, -29.60166, -10.2071,
  13.11834, 38.22106, 59.98977, 76.28748, 84.86707, 83.23065, 72.24286, 
    50.74245, 16.03397, -26.83344, -70.11647, -105.9174, -128.7831, 
    -137.0589, -132.006, -116.0477, -91.573, -65.9225, -40.8382, -13.82103,
  13.11821, 38.15613, 59.67234, 75.40578, 83.01276, 80.12503, 67.17565, 
    43.68682, 8.959417, -31.76498, -71.65201, -104.1217, -124.7371, 
    -132.2135, -127.6659, -113.1273, -90.5983, -66.00674, -41.00587, -13.91139,
  13.02355, 37.86329, 59.16221, 74.65988, 82.02097, 78.92241, 65.29362, 
    40.81419, 5.741602, -34.631, -73.57932, -104.7567, -124.1129, -130.7433, 
    -125.958, -111.7784, -90.0933, -65.93861, -40.92499, -13.88443,
  11.32619, 32.76077, 50.67513, 62.98497, 67.73914, 63.30512, 48.28465, 
    24.11987, -5.385161, -36.63582, -65.335, -87.8186, -102.0598, -107.7157, 
    -105.5208, -96.70057, -82.70698, -63.48643, -39.80992, -13.59205,
  11.14925, 32.24605, 49.86636, 61.95045, 66.58931, 62.22134, 47.65833, 
    24.35996, -4.084089, -34.27809, -62.27697, -84.66127, -99.36412, 
    -105.7874, -104.3717, -96.12457, -82.37784, -63.28226, -39.72206, 
    -13.56579,
  10.88813, 31.50476, 48.75818, 60.64318, 65.31243, 61.25799, 47.59411, 
    25.65779, -1.429946, -30.4262, -57.75721, -80.29189, -95.89642, 
    -103.5962, -103.3768, -95.88637, -82.23525, -63.11871, -39.66102, 
    -13.54348,
  10.50852, 30.43788, 47.19903, 58.87909, 63.71529, 60.23011, 47.90954, 
    27.82024, 2.349577, -25.38457, -52.1809, -75.20702, -92.19078, -101.6232, 
    -102.878, -96.15462, -82.30364, -62.9541, -39.58221, -13.50597,
  10.06445, 29.21246, 45.48198, 57.09265, 62.38165, 59.86744, 49.32035, 
    31.38589, 7.56664, -19.18434, -46.00835, -70.28177, -89.38877, -101.0308, 
    -103.8321, -97.59562, -83.08059, -63.09846, -39.59311, -13.4783,
  9.568386, 27.88424, 43.75979, 55.61941, 61.93172, 61.18333, 52.89923, 
    37.11209, 14.67563, -11.80515, -39.80424, -66.68553, -89.04987, 
    -103.3828, -107.4757, -101.0359, -85.22389, -63.92684, -39.74198, 
    -13.45525,
  7.81792, 22.81706, 35.87301, 45.66008, 51.01283, 51.30911, 46.0572, 
    34.12345, 17.32008, -2.352751, -23.36801, -44.26085, -62.3951, -74.53143, 
    -78.65536, -74.67769, -63.61718, -48.865, -31.25493, -10.69787,
  6.805508, 20.00689, 31.89069, 41.41726, 47.56139, 49.64371, 46.30203, 
    35.54575, 20.02802, 1.837487, -18.36294, -39.97929, -60.20417, -74.74669, 
    -80.81284, -78.22025, -67.93638, -52.16284, -32.88104, -11.15253,
  6.093643, 18.00475, 28.94953, 38.02238, 44.28236, 47.17881, 44.60117, 
    33.93987, 19.25903, 2.922509, -15.29974, -35.87211, -56.33062, -71.94724, 
    -79.44283, -78.56882, -70.21511, -54.02874, -33.405, -11.21848,
  5.829611, 17.26064, 27.83382, 36.64671, 42.75905, 45.77228, 43.03032, 
    31.60009, 17.02476, 2.116367, -14.03331, -32.86997, -52.56861, -68.42346, 
    -76.80151, -77.25057, -70.63613, -54.45082, -33.13451, -11.04475,
  6.047637, 17.91226, 28.90295, 38.09125, 44.52589, 47.87151, 45.07569, 
    32.86858, 17.53912, 2.317572, -13.79821, -32.60331, -52.49937, -68.66847, 
    -77.20267, -77.61071, -71.01836, -54.54338, -32.92459, -10.9314,
  6.713081, 19.86929, 32.05276, 42.3082, 49.67048, 53.72326, 51.34956, 
    38.88531, 22.04387, 4.258117, -14.81261, -36.30027, -57.94749, -74.44266, 
    -81.92529, -80.42073, -71.6759, -54.44554, -32.90019, -10.92455,
  7.683837, 22.70266, 36.54627, 48.18392, 56.5569, 60.99274, 58.7881, 
    46.16032, 27.28967, 5.654464, -17.92335, -43.1663, -66.64508, -82.67428, 
    -88.01162, -83.55855, -71.63493, -53.68177, -32.71988, -10.90888,
  8.739975, 25.74637, 41.2417, 54.03007, 62.8469, 66.67644, 63.646, 50.37846, 
    29.41883, 4.264261, -23.09889, -50.86705, -74.65926, -89.08847, 
    -91.94866, -84.8204, -70.15485, -51.98248, -32.0939, -10.77281,
  9.681756, 28.40042, 45.1342, 58.43813, 66.78931, 68.92625, 64.06192, 
    49.66174, 27.08981, -0.1233433, -29.19862, -57.21866, -79.50237, 
    -91.59099, -92.30421, -83.44069, -67.17006, -49.38908, -30.91271, 
    -10.45835,
  10.44449, 30.47625, 47.9287, 61.05053, 68.09114, 67.79978, 60.60421, 
    44.94398, 21.48207, -6.167258, -34.85173, -61.1735, -80.79659, -90.39958, 
    -89.52812, -79.84933, -63.08568, -46.14545, -29.22725, -9.96417,
  11.10049, 32.20081, 50.02696, 62.46287, 67.59078, 64.51591, 55.14739, 
    38.69369, 14.95468, -12.17204, -39.25092, -62.90253, -79.57539, 
    -86.98013, -85.01711, -75.01219, -58.19949, -42.28784, -27.09482, 
    -9.312143,
  12.24593, 35.56404, 55.43942, 69.72568, 76.32314, 73.19025, 62.29938, 
    44.12218, 16.53641, -17.43534, -53.49509, -86.18916, -109.8952, 
    -121.0378, -119.1875, -106.148, -84.36282, -60.93942, -37.78728, -12.78714,
  12.1894, 35.31118, 54.75244, 68.24779, 73.70975, 69.47481, 57.35146, 
    38.06198, 10.72504, -21.46257, -54.72911, -84.51211, -106.0839, -116.374, 
    -114.9116, -103.0873, -82.8949, -60.45173, -37.60901, -12.76061,
  12.08517, 34.97795, 54.13595, 67.28009, 72.35822, 67.85655, 55.24313, 
    35.33073, 7.96821, -23.69535, -56.08398, -84.81355, -105.3742, -114.9635, 
    -113.2945, -101.7633, -82.25846, -60.19827, -37.41318, -12.69423,
  10.31721, 29.69653, 45.47911, 55.68835, 58.79123, 53.96584, 40.9599, 
    21.7746, -0.478482, -23.91714, -46.47292, -65.91027, -80.16613, -87.8522, 
    -88.54669, -82.7382, -71.57464, -55.28088, -34.7856, -11.89308,
  10.17649, 29.29613, 44.88334, 55.00146, 58.15194, 53.51932, 40.92461, 
    22.29303, 0.5845557, -22.30959, -44.42626, -63.7086, -78.19817, 
    -86.43717, -87.79684, -82.53453, -71.62418, -55.41938, -34.93426, 
    -11.95102,
  10.00401, 28.82125, 44.22289, 54.32481, 57.65689, 53.37174, 41.42866, 
    23.60975, 2.593223, -19.65711, -41.3281, -60.63711, -75.75085, -85.04119, 
    -87.50409, -83.00961, -72.24805, -55.95029, -35.33583, -12.09095,
  9.769822, 28.17971, 43.33647, 53.41869, 56.98594, 53.14668, 42.03713, 
    25.267, 5.157599, -16.26168, -37.42085, -56.92556, -73.06812, -83.90104, 
    -87.84648, -84.25415, -73.49256, -56.86941, -35.9417, -12.28848,
  9.518674, 27.50361, 42.43499, 52.55614, 56.45486, 53.21637, 43.0213, 
    27.33452, 8.26611, -12.2259, -32.96323, -53.03261, -70.77567, -83.68593, 
    -89.38572, -86.66805, -75.75549, -58.4323, -36.7756, -12.53342,
  9.247168, 26.79553, 41.56298, 51.87661, 56.34913, 54.06169, 44.76764, 
    29.88778, 11.86094, -7.731082, -28.3421, -49.60862, -69.73389, -85.27313, 
    -92.77868, -90.59716, -79.27074, -60.67887, -37.68169, -12.74985,
  7.751707, 22.40922, 34.55101, 42.68325, 45.86968, 44.4355, 38.01484, 
    26.20829, 12.53616, -1.583939, -16.3831, -32.49581, -48.8551, -62.23698, 
    -69.19915, -68.18752, -59.5528, -45.85162, -29.08304, -9.930902,
  6.879671, 19.92398, 30.77422, 37.99081, 40.57122, 38.75914, 32.53825, 
    21.92595, 10.59617, -0.4079142, -12.48425, -27.33961, -44.3066, 
    -59.61491, -68.70809, -69.13889, -60.73371, -46.65014, -29.56649, 
    -10.07087,
  6.108829, 17.67609, 27.18354, 33.16532, 34.57904, 31.8262, 25.25449, 
    15.36563, 6.252826, -1.462493, -10.19717, -22.4716, -38.17311, -53.71679, 
    -64.16574, -66.41348, -59.59138, -45.88411, -28.8597, -9.785233,
  5.611314, 16.21311, 24.80033, 29.8531, 30.28969, 26.72161, 19.60714, 
    9.805275, 2.128082, -3.06076, -8.890978, -18.46454, -32.26522, -47.24408, 
    -58.48852, -62.45212, -57.73928, -44.75925, -27.84755, -9.392398,
  5.51461, 15.95713, 24.47193, 29.55619, 30.12288, 26.85922, 19.77632, 
    9.593904, 1.980536, -2.655878, -7.672947, -16.41883, -29.69073, 
    -44.69355, -56.46492, -61.27602, -57.72614, -44.92878, -27.66768, 
    -9.284822,
  5.873971, 17.06965, 26.45799, 32.63195, 34.53823, 32.74996, 26.47895, 
    15.73837, 6.725607, 0.2090493, -6.814336, -17.48575, -32.37779, -48.3056, 
    -60.03016, -64.07517, -59.73891, -46.23813, -28.3004, -9.46547,
  6.587636, 19.21301, 30.07795, 37.86345, 41.52748, 41.37921, 36.05052, 
    24.70897, 13.39714, 3.444856, -7.364823, -21.60771, -39.17494, -56.03173, 
    -66.70327, -68.47221, -61.74116, -47.19577, -28.90537, -9.668678,
  7.421476, 21.65831, 34.01518, 43.17326, 48.03525, 48.60886, 43.59113, 
    31.70932, 18.14742, 4.74961, -9.837425, -27.43822, -47.03008, -63.77882, 
    -72.42738, -71.32551, -61.79665, -46.59824, -28.74041, -9.649698,
  8.13949, 23.69206, 37.05672, 46.81262, 51.7748, 51.78103, 46.25223, 
    34.03352, 19.02108, 3.340354, -13.70875, -33.15806, -53.11211, -68.44971, 
    -74.67579, -71.10484, -59.43036, -44.26813, -27.58212, -9.316737,
  8.647326, 25.03999, 38.77496, 48.25884, 52.2733, 50.79487, 44.35684, 
    32.14115, 16.61147, 0.0007258654, -17.91875, -37.45145, -56.15863, 
    -69.26733, -73.28461, -68.10631, -55.32094, -40.74105, -25.61485, 
    -8.706841,
  9.006442, 25.89411, 39.51223, 48.04538, 50.37455, 47.05519, 39.99961, 
    28.44907, 13.03952, -3.842398, -21.75689, -40.25426, -56.77903, 
    -67.39057, -69.54239, -63.31309, -49.89931, -36.16757, -22.93051, 
    -7.848431,
  9.923043, 28.57387, 43.76311, 53.51848, 56.253, 50.95401, 41.22508, 
    29.45079, 13.98842, -4.78276, -26.84653, -50.88745, -73.0285, -88.11611, 
    -92.63306, -86.19309, -70.51862, -51.85058, -32.41204, -10.99852,
  9.731216, 27.89881, 42.33522, 51.00462, 52.52843, 46.53993, 36.69537, 
    24.96459, 9.995129, -7.584741, -27.82951, -49.7501, -70.01787, -84.05702, 
    -88.56583, -82.85751, -68.15121, -50.3562, -31.63807, -10.77402,
  9.577699, 27.4039, 41.40807, 49.54416, 50.53785, 44.31149, 34.34259, 
    22.50776, 7.845851, -9.076052, -28.50839, -49.6229, -69.18856, -82.73737, 
    -87.07923, -81.54398, -67.2677, -49.77962, -31.24887, -10.64287,
  8.839197, 25.28971, 38.26797, 46.03637, 47.53398, 42.61305, 31.73162, 
    17.06872, 1.114877, -15.40588, -31.95193, -47.57612, -60.70152, 
    -69.51564, -72.68675, -69.85309, -61.63387, -48.21758, -30.57294, 
    -10.48969,
  8.75405, 25.05899, 37.96505, 45.77573, 47.44525, 42.78025, 32.22663, 
    17.85725, 2.072512, -14.2912, -30.65958, -46.18004, -59.41294, -68.59213, 
    -72.28067, -69.91815, -61.92865, -48.56541, -30.85912, -10.59555,
  8.686446, 24.8955, 37.81225, 45.77832, 47.74103, 43.41708, 33.28771, 
    19.29728, 3.706628, -12.46027, -28.64002, -44.18889, -57.86034, 
    -67.86449, -72.50235, -70.85321, -63.03012, -49.52005, -31.53148, 
    -10.82879,
  8.601249, 24.68853, 37.60818, 45.73309, 47.99488, 44.02039, 34.33574, 
    20.78493, 5.523359, -10.25208, -26.0946, -41.71336, -56.10956, -67.37122, 
    -73.35059, -72.61458, -64.91943, -51.0406, -32.50272, -11.14994,
  8.526059, 24.51627, 37.4663, 45.76512, 48.32607, 44.74467, 35.42004, 
    22.19016, 7.378747, -7.818807, -23.23857, -39.05788, -54.52459, 
    -67.45995, -75.07439, -75.35157, -67.8358, -53.2785, -33.71837, -11.52028,
  8.435903, 24.31505, 37.31572, 45.84048, 48.77357, 45.72738, 36.57351, 
    23.34503, 9.076443, -5.402591, -20.44394, -36.74083, -53.68666, 
    -68.62466, -77.92943, -79.04592, -71.66289, -56.02236, -34.91367, 
    -11.83086,
  7.116107, 20.41097, 30.97964, 37.39895, 39.085, 37.0207, 30.84752, 
    20.28575, 9.179472, -1.460941, -12.33617, -24.66185, -38.32754, 
    -50.96646, -59.05473, -60.12631, -53.60585, -41.40252, -26.17973, 
    -8.940233,
  6.328864, 18.116, 27.31287, 32.45525, 32.85389, 29.45442, 22.97036, 
    13.94504, 5.483255, -1.979022, -10.04084, -20.57153, -33.80259, 
    -47.27214, -56.7856, -58.94976, -52.37472, -40.32126, -25.72815, -8.804177,
  5.515957, 15.69007, 23.26743, 26.71801, 25.35775, 20.40128, 13.50645, 
    5.899839, 0.1632862, -3.926353, -8.721521, -16.47745, -27.76881, 
    -40.55719, -50.7153, -54.3138, -49.02446, -37.83603, -24.17405, -8.268291,
  4.871851, 13.75775, 20.01749, 22.07, 19.27456, 13.18992, 5.973952, 
    -0.7217875, -4.355925, -5.654787, -7.512819, -12.46441, -21.48012, 
    -33.15081, -43.70642, -48.93073, -45.77057, -35.71378, -22.69754, 
    -7.742294,
  4.575942, 12.90453, 18.69827, 20.41041, 17.43839, 11.49559, 4.470429, 
    -2.008194, -4.863231, -5.01441, -5.607974, -9.348392, -17.49501, 
    -29.01445, -40.26373, -46.82179, -45.39542, -35.85085, -22.56682, 
    -7.661644,
  4.731189, 13.43566, 19.80965, 22.42648, 20.70019, 16.22211, 9.957082, 
    3.022661, -0.6350729, -1.756277, -3.397413, -8.279629, -17.69004, 
    -30.42495, -42.4958, -49.37904, -48.21157, -38.12281, -23.74857, -8.019545,
  5.262783, 15.08377, 22.76027, 26.99603, 27.18566, 24.60768, 19.21207, 
    11.36566, 5.766035, 2.190887, -2.061441, -9.653921, -21.67579, -36.2313, 
    -48.62169, -54.45908, -51.89733, -40.63306, -25.1576, -8.467821,
  5.938138, 17.11032, 26.17804, 31.91177, 33.65544, 32.3476, 27.43726, 
    18.69741, 10.96969, 4.678428, -2.436179, -12.94267, -27.53269, -43.33488, 
    -54.99886, -58.67273, -53.73712, -41.46207, -25.68626, -8.650285,
  6.505249, 18.74404, 28.72448, 35.19942, 37.47308, 36.29318, 31.36084, 
    22.22584, 13.05748, 4.785314, -4.465725, -17.04639, -33.05212, -48.75013, 
    -58.67304, -59.83967, -52.56206, -39.9347, -24.87965, -8.40958,
  6.848775, 19.64409, 29.84926, 36.14227, 37.8807, 35.94173, 30.81118, 
    21.96855, 12.28581, 2.987184, -7.419206, -20.84285, -36.73491, -51.01275, 
    -58.74054, -57.8126, -48.9274, -36.57888, -22.92569, -7.786311,
  7.014023, 19.95085, 29.80324, 35.14893, 35.58339, 32.55247, 27.62355, 
    19.9202, 10.38202, 0.4630113, -10.64862, -24.04996, -38.64719, -50.645, 
    -56.06594, -53.44194, -43.37341, -31.66743, -19.95868, -6.819208,
  7.775893, 22.16751, 33.26448, 39.40639, 39.56662, 33.5242, 25.51431, 
    18.49062, 10.90303, 1.875054, -10.33834, -26.64912, -45.23282, -61.44515, 
    -70.32628, -69.44512, -59.24542, -44.76016, -28.3478, -9.669513,
  7.474876, 21.16634, 31.31479, 36.26618, 35.31968, 28.92825, 21.44702, 
    15.05514, 7.994452, -0.2444854, -11.27049, -26.06388, -43.07274, 
    -58.1185, -66.59531, -65.95711, -56.18499, -42.47834, -27.11323, -9.293643,
  7.270782, 20.51418, 30.11576, 34.43565, 32.93575, 26.40609, 19.0712, 
    12.86288, 6.203241, -1.412897, -11.70823, -25.80004, -42.22947, 
    -56.87988, -65.19827, -64.6362, -55.10042, -41.64848, -26.57652, -9.114077,
  6.834525, 19.36126, 28.73261, 33.60782, 33.51431, 28.93327, 20.76395, 
    11.0641, 1.644319, -7.684289, -17.56132, -28.26898, -39.0858, -48.28066, 
    -53.84572, -54.43816, -49.86035, -39.99621, -25.74092, -8.894349,
  6.823623, 19.35478, 28.80471, 33.86026, 34.02966, 29.70218, 21.71646, 
    12.04642, 2.487047, -6.992157, -16.93401, -27.64454, -38.51132, 
    -47.90304, -53.80617, -54.74951, -50.35189, -40.49935, -26.12184, 
    -9.032221,
  6.881206, 19.55897, 29.23532, 34.60565, 35.12848, 31.06519, 23.22801, 
    13.52201, 3.742407, -5.90639, -15.90334, -26.69339, -37.8581, -47.83718, 
    -54.4803, -56.02939, -51.79972, -41.75828, -26.97797, -9.327402,
  6.957781, 19.82006, 29.75192, 35.43866, 36.27959, 32.42836, 24.64512, 
    14.82497, 4.873235, -4.795547, -14.68119, -25.49352, -37.0914, -47.9567, 
    -55.67236, -58.05326, -54.05946, -43.64708, -28.15922, -9.718292,
  7.054007, 20.13667, 30.34138, 36.32445, 37.43397, 33.80405, 25.92216, 
    15.78046, 5.723088, -3.818997, -13.48803, -24.3152, -36.45224, -48.38866, 
    -57.36153, -60.7195, -57.17429, -46.18783, -29.53973, -10.14269,
  7.117373, 20.36448, 30.8052, 37.06249, 38.42747, 35.07262, 26.88566, 
    16.16025, 6.102433, -3.209362, -12.70124, -23.65713, -36.40997, 
    -49.39657, -59.50219, -63.70565, -60.7122, -48.96496, -30.8043, -10.48227,
  5.923339, 16.81493, 25.0105, 29.35151, 29.74521, 27.71693, 22.78291, 
    14.43784, 6.21698, -1.222079, -8.633402, -17.25327, -27.53007, -38.15732, 
    -46.28081, -49.05508, -44.87309, -34.82441, -21.99065, -7.523679,
  5.164903, 14.56263, 21.28683, 24.11183, 22.85565, 19.02291, 13.71314, 
    7.288527, 1.663842, -3.062102, -8.12555, -14.92231, -24.00348, -34.21495, 
    -42.60667, -45.77587, -41.23585, -31.87014, -20.56862, -7.092727,
  4.276338, 11.87682, 16.72595, 17.56284, 14.30154, 8.761534, 3.295933, 
    -1.162295, -3.962855, -5.64027, -7.856315, -12.04011, -18.84507, 
    -27.56433, -35.66737, -39.58099, -35.91804, -27.80364, -18.19961, 
    -6.309705,
  3.484886, 9.478548, 12.6466, 11.72681, 6.79357, 0.08733654, -5.338189, 
    -8.239074, -8.572546, -7.418808, -6.815553, -8.284842, -12.70561, 
    -19.9307, -27.94902, -33.14272, -31.41755, -24.72784, -16.26566, -5.650873,
  3.016053, 8.09356, 10.41039, 8.762714, 3.335524, -3.39202, -8.434045, 
    -10.51381, -9.425457, -6.594359, -4.33655, -4.321223, -7.677429, 
    -14.63836, -23.4113, -30.21234, -30.55335, -24.67815, -16.1256, -5.584209,
  3.004693, 8.129995, 10.70629, 9.638168, 5.122486, -0.4235725, -4.807576, 
    -6.996292, -5.931987, -3.10057, -0.9520967, -1.326776, -5.533747, 
    -13.82026, -24.11265, -32.27456, -33.85085, -27.70169, -17.8129, -6.118705,
  3.389602, 9.36449, 13.03441, 13.41532, 10.63268, 6.817643, 3.04094, 
    -0.08724689, -0.2834868, 1.244965, 2.03393, -0.02584505, -6.404163, 
    -16.98966, -28.92219, -37.60086, -39.08235, -31.80871, -20.13287, -6.86014,
  3.937701, 11.05343, 16.01422, 17.90968, 16.77013, 14.38987, 10.95069, 
    6.619894, 4.676962, 4.454074, 3.540095, -0.5423121, -9.382366, -22.18837, 
    -35.02328, -42.97896, -43.06645, -34.5147, -21.64828, -7.344712,
  4.385313, 12.38277, 18.21693, 21.00486, 20.72985, 18.97637, 15.6612, 
    10.61245, 7.289676, 5.603189, 3.247169, -2.533962, -13.23896, -27.21765, 
    -39.64475, -45.78612, -43.77255, -34.42341, -21.5495, -7.310402,
  4.597722, 12.94554, 18.95965, 21.76245, 21.42234, 19.59887, 16.50311, 
    11.61654, 7.661972, 5.000222, 1.567207, -5.327989, -16.79072, -30.46051, 
    -41.29003, -45.21275, -41.21948, -31.72811, -19.87657, -6.758083,
  4.598682, 12.81136, 18.35984, 20.38578, 19.26363, 17.09644, 14.74345, 
    11.05214, 7.106138, 3.602674, -0.9369373, -8.564102, -19.71003, 
    -31.73058, -40.12498, -41.72113, -35.89076, -26.72325, -16.75768, 
    -5.723197,
  5.220697, 14.61185, 21.1166, 23.56418, 21.59103, 15.67735, 10.06494, 
    7.738679, 7.270211, 6.93301, 4.006122, -3.922294, -17.10199, -32.47034, 
    -44.81197, -49.83552, -46.11019, -36.68332, -23.80652, -8.202357,
  4.809438, 13.29559, 18.71043, 19.97044, 17.0991, 11.12782, 6.528215, 
    5.284596, 5.319762, 5.408968, 3.10075, -3.930511, -15.96378, -30.16871, 
    -41.68585, -46.32091, -42.32216, -33.51794, -22.05329, -7.656395,
  4.544848, 12.46265, 17.22392, 17.7982, 14.41838, 8.435273, 4.226945, 
    3.399753, 3.857809, 4.467124, 2.76079, -3.675175, -15.20964, -29.0657, 
    -40.40046, -44.98948, -41.00278, -32.39314, -21.3476, -7.421937,
  3.102924, 8.457497, 11.61709, 12.08376, 10.25831, 7.166918, 3.708705, 
    1.328269, 0.9323757, 1.526361, 1.477033, -0.8314247, -6.157395, 
    -13.77406, -21.6013, -27.17801, -28.80285, -25.33205, -17.17676, -6.082424,
  3.222309, 8.835775, 12.29975, 13.09855, 11.55966, 8.597154, 5.054698, 
    2.381084, 1.560628, 1.740963, 1.379617, -1.112887, -6.518537, -14.17565, 
    -22.07363, -27.75652, -29.43324, -25.90284, -17.57342, -6.221776,
  3.465415, 9.573509, 13.53727, 14.79078, 13.56691, 10.66433, 6.877778, 
    3.7021, 2.275124, 1.942951, 1.24829, -1.446166, -7.032276, -14.94544, 
    -23.19124, -29.20578, -31.00066, -27.25524, -18.45145, -6.51995,
  3.747937, 10.42019, 14.92224, 16.62008, 15.65707, 12.76291, 8.590712, 
    4.734761, 2.641761, 1.80968, 0.8422251, -1.977514, -7.697871, -15.89287, 
    -24.58766, -31.07508, -33.15133, -29.10917, -19.56592, -6.884126,
  4.023936, 11.24574, 16.26382, 18.37611, 17.66268, 14.87092, 10.22061, 
    5.462448, 2.657363, 1.273978, -0.04256058, -3.007006, -8.766567, 
    -17.07189, -26.07747, -33.05696, -35.70704, -31.34672, -20.75589, 
    -7.246078,
  4.208562, 11.81713, 17.23932, 19.71872, 19.26562, 16.65731, 11.46235, 
    5.694386, 2.201909, 0.1574985, -1.741838, -4.988793, -10.63573, 
    -18.61628, -27.42592, -34.61145, -37.9701, -33.42424, -21.76031, -7.522312,
  3.084622, 8.50541, 11.9599, 13.02502, 12.35377, 11.73754, 10.20825, 
    6.488666, 2.9283, -0.1357715, -3.162027, -6.900344, -11.92404, -18.09862, 
    -24.17034, -27.96963, -27.00541, -21.07063, -13.24519, -4.562394,
  2.263031, 6.063285, 7.935726, 7.423015, 5.085873, 2.598532, 0.9549894, 
    -0.5069747, -1.92396, -3.257894, -4.902785, -7.231209, -10.56737, 
    -14.94188, -19.51151, -22.28584, -20.30361, -15.63344, -10.47477, 
    -3.709837,
  1.20703, 2.894368, 2.660997, 0.1122646, -4.055573, -8.003352, -9.37543, 
    -8.552591, -7.479248, -6.486534, -6.009843, -6.16496, -7.162142, 
    -9.344538, -12.42518, -14.70425, -12.74797, -9.597946, -7.01826, -2.583498,
  0.1939453, -0.1555083, -2.428426, -6.913058, -12.67782, -17.56586, 
    -18.48123, -15.67177, -12.06141, -8.409945, -5.369192, -3.048186, 
    -1.75358, -2.206123, -4.594156, -7.402463, -6.764389, -5.216641, 
    -4.401246, -1.715911,
  -0.4939173, -2.208097, -5.787043, -11.40045, -17.9207, -22.94131, 
    -23.24932, -19.02679, -13.4085, -7.574806, -2.49805, 1.537425, 4.020732, 
    3.945572, 0.9153719, -3.473344, -4.939955, -4.547572, -4.045265, -1.605728,
  -0.689423, -2.753081, -6.54715, -12.14092, -18.32863, -22.63891, -22.34797, 
    -17.61874, -11.03822, -4.089127, 1.91921, 6.400752, 8.582792, 7.323348, 
    2.345404, -4.354152, -8.095992, -7.991531, -6.181767, -2.32405,
  -0.4469835, -1.9709, -5.064682, -9.737239, -14.82151, -17.94494, -17.32068, 
    -13.13261, -6.724959, 0.3553798, 6.475446, 10.57091, 11.46702, 7.974159, 
    0.2578812, -8.946599, -14.59705, -13.90558, -9.719993, -3.49098,
  -0.00469172, -0.5964935, -2.622926, -6.066508, -9.851243, -11.76627, 
    -11.11067, -8.164885, -2.698179, 3.962851, 9.896619, 13.38525, 12.70136, 
    6.687685, -3.730877, -14.83116, -21.41347, -19.57532, -12.97614, -4.543003,
  0.3597245, 0.5235062, -0.6646309, -3.166719, -5.963084, -6.948813, 
    -6.305117, -4.54079, -0.170002, 5.897066, 11.54847, 14.41583, 12.26963, 
    4.173683, -7.972095, -19.54586, -25.65004, -22.60767, -14.56419, -5.032651,
  0.4825237, 0.8899727, -0.03475046, -2.199472, -4.514563, -4.824447, 
    -3.846178, -2.538145, 1.036363, 6.420363, 11.51766, 13.60599, 10.29887, 
    1.132699, -11.13193, -21.54518, -25.98895, -22.0987, -13.98374, -4.80192,
  0.3431102, 0.4280353, -0.8827662, -3.366275, -5.665191, -5.41691, 
    -3.445662, -1.444644, 1.826777, 6.293154, 10.21047, 11.09827, 6.992207, 
    -1.920255, -12.51173, -20.30033, -22.12159, -17.82017, -11.08517, -3.80191,
  0.8190162, 1.794657, 1.128005, -1.375637, -5.180418, -9.226459, -10.52838, 
    -6.638632, 1.60778, 11.7855, 20.6669, 24.82508, 21.78456, 11.55963, 
    -2.546485, -15.29263, -22.32898, -22.07819, -15.65949, -5.591683,
  0.2741131, 0.1293259, -1.68127, -5.180151, -9.515566, -13.46721, -13.39091, 
    -7.919937, 0.8080113, 11.04257, 19.91557, 24.15514, 21.45861, 12.01296, 
    -0.8981438, -12.21555, -17.58732, -17.49771, -13.05243, -4.762638,
  -0.088094, -0.9763546, -3.543673, -7.701731, -12.3931, -16.23121, 
    -15.51883, -9.361833, -0.2234296, 10.35535, 19.60048, 24.22974, 21.89646, 
    12.76039, 0.1190853, -10.90683, -15.86657, -15.84417, -12.04867, -4.432335,
  0.3540901, 0.5430806, -0.4588141, -2.52788, -4.872553, -6.478677, 
    -6.804512, -4.902308, -0.2818677, 5.833588, 11.55776, 14.79416, 13.98749, 
    8.93501, 1.114565, -6.88088, -12.54024, -13.77856, -10.36278, -3.83884,
  0.5581169, 1.162525, 0.5784025, -1.120711, -3.229258, -4.816748, -5.369473, 
    -3.888097, 0.2239228, 5.847315, 11.16175, 14.10817, 13.15767, 8.100473, 
    0.3528852, -7.565419, -13.15295, -14.2708, -10.67283, -3.943034,
  0.8931487, 2.155417, 2.173759, 0.9435239, -0.9217944, -2.560665, -3.513936, 
    -2.692909, 0.6988135, 5.680714, 10.51258, 13.14564, 12.02507, 6.886483, 
    -0.9237528, -8.913204, -14.52101, -15.41511, -11.37443, -4.175041,
  1.25343, 3.216796, 3.858963, 3.090365, 1.445461, -0.238019, -1.694801, 
    -1.716309, 0.8489504, 5.103343, 9.397356, 11.72502, 10.51423, 5.40799, 
    -2.384089, -10.45689, -16.23476, -16.88333, -12.20353, -4.437334,
  1.573975, 4.169664, 5.394819, 5.090395, 3.732536, 2.184141, 0.2085886, 
    -0.8467991, 0.7814673, 4.132207, 7.672402, 9.575583, 8.363124, 3.567511, 
    -3.894337, -11.92316, -18.09526, -18.55733, -13.04886, -4.684556,
  1.768693, 4.780705, 6.464298, 6.60839, 5.602054, 4.293192, 1.813046, 
    -0.3063078, 0.3484629, 2.583755, 5.046513, 6.332521, 5.271003, 1.298713, 
    -5.188128, -12.75691, -19.37487, -19.92174, -13.74504, -4.878076,
  0.6459655, 1.529908, 1.467807, 0.6304374, -0.04680729, 0.9433541, 2.207302, 
    1.91543, 1.483652, 1.158858, 0.7026135, -0.2769339, -2.183773, -5.223254, 
    -9.025831, -12.33278, -12.81289, -9.764692, -5.935518, -2.060142,
  -0.2399365, -1.06752, -2.706618, -5.016067, -7.214762, -8.000151, 
    -6.699634, -4.700749, -3.309388, -2.40726, -1.97241, -1.853033, 
    -2.064579, -2.879396, -4.387143, -5.801524, -4.723313, -3.088355, 
    -2.450922, -0.9773222,
  -1.396388, -4.48447, -8.233901, -12.41538, -16.19082, -18.25247, -16.55145, 
    -12.30806, -8.735569, -5.915996, -3.731402, -1.705757, 0.3132973, 
    1.835843, 2.287981, 2.062168, 3.735967, 3.89157, 1.577443, 0.3395922,
  -2.530578, -7.851238, -13.70723, -19.72804, -24.89652, -27.73653, 
    -25.47244, -19.24059, -13.28525, -8.010055, -3.449069, 0.890857, 
    5.091816, 8.37687, 9.793737, 9.524288, 10.39825, 9.001542, 4.621746, 
    1.347128,
  -3.338535, -10.24516, -17.56908, -24.78933, -30.70237, -33.66225, 
    -30.72876, -22.95642, -14.90811, -7.37753, -0.7130988, 5.388696, 
    10.82288, 14.58491, 15.55255, 13.94862, 12.94623, 10.27767, 5.273367, 
    1.541493,
  -3.636559, -11.11225, -18.89887, -26.35357, -32.1518, -34.56921, -31.0318, 
    -22.49892, -13.16328, -4.163721, 3.780598, 10.64815, 16.07067, 18.8919, 
    18.02763, 14.0026, 10.451, 7.118241, 3.156121, 0.799728,
  -3.469657, -10.59344, -17.95651, -24.84659, -29.89798, -31.39002, 
    -27.56084, -19.26877, -9.627779, 0.04735076, 8.656704, 15.6859, 20.34008, 
    21.28828, 17.63698, 10.48702, 4.089684, 0.7712936, -0.8401685, -0.5558819,
  -3.068513, -9.37964, -15.89004, -21.86225, -25.93583, -26.41297, -22.63393, 
    -15.41469, -6.257339, 3.580536, 12.63706, 19.73575, 23.46058, 22.24222, 
    15.52431, 5.255746, -3.633527, -6.32973, -5.095848, -1.963056,
  -2.710012, -8.294256, -14.04284, -19.20248, -22.40621, -21.928, -18.26791, 
    -12.36126, -4.048501, 5.661137, 15.02237, 22.16374, 25.01255, 21.82862, 
    12.59304, 0.2396412, -9.880211, -11.54767, -7.989837, -2.882885,
  -2.573944, -7.873605, -13.28644, -18.00265, -20.56626, -19.1308, -15.24069, 
    -10.21636, -2.717169, 6.571482, 15.79855, 22.61011, 24.52996, 19.9263, 
    9.48905, -3.086301, -12.63767, -13.18725, -8.566754, -3.01184,
  -2.719024, -8.305286, -13.94702, -18.68718, -20.85807, -18.47694, 
    -13.70217, -8.500858, -1.463992, 7.018227, 15.2808, 20.98427, 21.80668, 
    16.64391, 6.873076, -3.672591, -10.66212, -10.22407, -6.251934, -2.16908,
  -2.281462, -7.0655, -12.20684, -17.2247, -21.2347, -23.18304, -21.58496, 
    -14.44648, -1.858271, 13.54568, 28.53704, 39.5726, 43.45561, 38.54998, 
    26.08185, 10.26708, -3.587853, -10.16928, -8.912739, -3.422637,
  -2.871952, -8.823112, -15.03977, -20.86868, -25.24942, -27.25156, -24.2519, 
    -15.2694, -2.138092, 13.25209, 28.04042, 38.80945, 42.54102, 37.93935, 
    26.55178, 12.65501, 1.486844, -4.751794, -5.766737, -2.408675,
  -3.293231, -10.07851, -17.0668, -23.48077, -28.11678, -30.0264, -26.32709, 
    -16.50764, -2.954001, 12.71202, 27.75837, 38.78325, 42.75782, 38.40245, 
    27.32304, 13.89213, 3.473377, -2.708988, -4.547235, -2.009413,
  -2.367146, -7.185934, -11.96378, -16.02367, -18.42569, -18.42423, 
    -15.96508, -10.5317, -1.882942, 8.687696, 19.24405, 27.48224, 31.32948, 
    29.74384, 23.31363, 14.1851, 5.185902, -0.7323136, -2.492104, -1.220699,
  -2.094337, -6.378994, -10.67392, -14.37089, -16.6017, -16.6581, -14.49718, 
    -9.533908, -1.416988, 8.623186, 18.69746, 26.54804, 30.16572, 28.55793, 
    22.2896, 13.40493, 4.623744, -1.090333, -2.663582, -1.268959,
  -1.712175, -5.262472, -8.924524, -12.17453, -14.21278, -14.3516, -12.62659, 
    -8.360488, -0.9931019, 8.322847, 17.77504, 25.1699, 28.55751, 26.96109, 
    20.87272, 12.20293, 3.565586, -1.887637, -3.08119, -1.394581,
  -1.333383, -4.153355, -7.180429, -9.971118, -11.78494, -11.92836, 
    -10.68553, -7.276004, -0.7861682, 7.651948, 16.3311, 23.19229, 26.39943, 
    24.98225, 19.27719, 10.93734, 2.359096, -2.840142, -3.52661, -1.5178,
  -1.020464, -3.215413, -5.644728, -7.926018, -9.379623, -9.304094, 
    -8.509622, -6.112633, -0.645497, 6.677169, 14.29366, 20.42399, 23.47653, 
    22.50235, 17.54527, 9.760921, 1.128705, -3.905934, -3.989862, -1.634844,
  -0.8415418, -2.631714, -4.567196, -6.322046, -7.333634, -6.966979, 
    -6.587178, -5.192536, -0.8146189, 5.162647, 11.39453, 16.59377, 19.60898, 
    19.54827, 15.98004, 9.221197, 0.5745964, -4.634977, -4.402159, -1.752501,
  -1.949086, -5.770803, -9.191841, -11.51109, -11.77782, -9.038924, 
    -5.051541, -2.052301, 0.5039978, 2.811693, 4.764043, 6.217022, 6.964818, 
    6.725241, 5.336802, 3.200819, 2.030707, 2.46991, 2.152764, 0.7491895,
  -2.863394, -8.414327, -13.34704, -17.02068, -18.70837, -17.69312, 
    -13.61256, -8.378898, -4.21207, -0.9436412, 1.637795, 3.96905, 6.295942, 
    8.375849, 9.66788, 10.01146, 10.87462, 9.925072, 6.116828, 1.990631,
  -4.063072, -11.9056, -18.85403, -24.20447, -27.27849, -27.46498, -22.98283, 
    -15.62502, -9.530056, -4.61795, -0.5282133, 3.505924, 7.914355, 12.31209, 
    15.77893, 17.77467, 19.76047, 17.48555, 10.53065, 3.443344,
  -5.261659, -15.41066, -24.40928, -31.42382, -35.69337, -36.56834, -31.5273, 
    -22.29412, -14.04003, -6.908944, -0.6408556, 5.551507, 12.0358, 18.1954, 
    22.81335, 25.16235, 26.84212, 23.15281, 13.93396, 4.575633,
  -6.151675, -18.01248, -28.50983, -36.65652, -41.56484, -42.52054, 
    -36.81643, -26.08719, -15.86324, -6.606111, 1.679017, 9.603236, 17.35988, 
    24.13539, 28.5656, 29.93323, 30.09677, 25.12023, 14.97877, 4.894926,
  -6.539654, -19.13829, -30.23222, -38.69492, -43.52576, -43.98729, -37.689, 
    -26.13929, -14.59905, -3.841373, 5.797343, 14.62842, 22.60082, 28.74707, 
    31.68246, 30.87236, 28.56615, 22.65704, 13.17207, 4.231703,
  -6.455844, -18.88517, -29.76599, -37.87273, -42.1186, -41.76538, -35.1759, 
    -23.70464, -11.67392, -0.05632466, 10.45687, 19.73018, 27.31859, 
    32.03815, 32.52677, 28.58952, 23.05466, 16.62122, 9.160913, 2.828672,
  -6.109169, -17.86867, -28.10987, -35.54839, -39.01982, -37.74909, 
    -31.21417, -20.65501, -8.845101, 3.210856, 14.46597, 24.18523, 31.3371, 
    34.39211, 32.01264, 24.50527, 15.45482, 8.957361, 4.339704, 1.189644,
  -5.757949, -16.83935, -26.44304, -33.24102, -35.96914, -33.72851, -27.3595, 
    -18.13708, -6.969859, 5.244459, 17.14639, 27.34651, 34.14573, 35.63802, 
    30.59357, 19.9798, 8.112643, 2.104271, 0.3401742, -0.1193147,
  -5.584229, -16.32217, -25.56849, -31.92173, -33.96343, -30.58447, 
    -24.10282, -16.08183, -5.688425, 6.340563, 18.45494, 28.74331, 34.99199, 
    35.11943, 28.24034, 16.04786, 3.184401, -1.793131, -1.533637, -0.6678361,
  -5.682883, -16.59732, -25.92166, -32.1071, -33.54179, -28.96494, -21.79416, 
    -14.09952, -4.245836, 7.173169, 18.64496, 28.11362, 33.29689, 32.38958, 
    25.15835, 13.84925, 2.742268, -0.8033042, -0.1734149, -0.09994853,
  -5.245359, -15.39442, -24.36321, -31.10114, -34.63809, -34.18164, 
    -29.99632, -20.47152, -4.751597, 14.46218, 34.05703, 50.6081, 60.68818, 
    61.6332, 52.729, 36.2345, 17.00712, 3.709948, -0.7762089, -0.7700984,
  -5.839402, -17.1264, -27.0625, -34.46764, -38.35255, -38.2567, -32.77014, 
    -21.17838, -4.762419, 14.53307, 33.9436, 50.11283, 59.72166, 60.47383, 
    52.23982, 37.75371, 22.02578, 9.664068, 2.761512, 0.3885734,
  -6.306665, -18.48647, -29.17505, -37.08442, -41.17278, -41.10068, 
    -34.91881, -22.34789, -5.455878, 14.12023, 33.7542, 50.10423, 59.8495, 
    60.7471, 52.79216, 38.88816, 24.23817, 12.07881, 4.180893, 0.8514097,
  -4.832011, -14.09408, -22.00958, -27.48769, -29.65515, -28.16708, 
    -23.46111, -15.3374, -3.665905, 10.27948, 24.62882, 37.06224, 45.26057, 
    47.58131, 43.70614, 34.92226, 23.75043, 13.62674, 6.475022, 1.813102,
  -4.515366, -13.175, -20.58687, -25.7285, -27.76815, -26.35659, -21.9459, 
    -14.27651, -3.118451, 10.2829, 24.09298, 36.04558, 43.90881, 46.13239, 
    42.42551, 33.98855, 23.17207, 13.36167, 6.426697, 1.818275,
  -4.132635, -12.06375, -18.8621, -23.57824, -25.4234, -24.04021, -19.99886, 
    -12.97074, -2.529037, 10.10721, 23.1757, 34.51328, 42.01569, 44.2246, 
    40.81978, 32.82602, 22.34943, 12.88779, 6.293097, 1.802844,
  -3.781997, -11.0327, -17.22576, -21.47717, -23.04657, -21.5658, -17.89474, 
    -11.6333, -2.031428, 9.665478, 21.7963, 32.3807, 39.51846, 41.8626, 
    38.99725, 31.63272, 21.48367, 12.36149, 6.184777, 1.806738,
  -3.501496, -10.17574, -15.779, -19.48296, -20.62021, -18.84171, -15.50122, 
    -10.12854, -1.510421, 9.017149, 19.92717, 29.54267, 36.28683, 38.95661, 
    36.94455, 30.44378, 20.59505, 11.71707, 5.990633, 1.783798,
  -3.329994, -9.600215, -14.68348, -17.82265, -18.48939, -16.42679, 
    -13.41454, -8.906501, -1.332992, 7.846396, 17.2912, 25.78785, 32.23796, 
    35.62341, 35.01597, 29.81635, 20.35279, 11.35442, 5.723616, 1.697734,
  -4.373226, -12.50062, -18.79894, -22.18613, -21.90207, -17.62812, -11.3231, 
    -5.420469, -0.1307018, 4.672447, 8.902981, 12.52906, 15.49052, 17.55889, 
    18.34944, 17.65946, 16.42173, 14.71521, 10.44105, 3.67592,
  -5.253238, -15.03104, -22.75634, -27.44853, -28.59292, -26.06107, 
    -19.67798, -11.62584, -4.811531, 0.9032734, 5.714192, 10.12062, 14.51711, 
    18.79867, 22.32251, 24.36398, 25.43979, 22.45778, 14.60808, 4.985455,
  -6.417472, -18.39049, -27.9925, -34.22537, -36.69028, -35.39622, -28.68377, 
    -18.63226, -10.05285, -2.837034, 3.357617, 9.330964, 15.65911, 22.15175, 
    27.88275, 31.80786, 34.35452, 30.22656, 19.18387, 6.500534,
  -7.603059, -21.82097, -33.34007, -41.06755, -44.60139, -43.98679, -36.7827, 
    -25.00715, -14.5045, -5.311388, 2.858932, 10.83612, 19.14132, 27.38576, 
    34.3983, 38.97566, 41.62457, 36.25013, 22.83751, 7.725064,
  -8.514031, -24.44714, -37.38456, -46.10277, -50.14674, -49.58628, 
    -41.77833, -28.65839, -16.44283, -5.395427, 4.585005, 14.19385, 23.79645, 
    32.81824, 39.94118, 43.93936, 45.49933, 38.91164, 24.32488, 8.195486,
  -8.957323, -25.70613, -39.24146, -48.20866, -52.0949, -51.02972, -42.6785, 
    -28.8455, -15.51386, -3.181495, 8.009516, 18.51733, 28.49613, 37.21799, 
    43.29944, 45.59097, 45.04453, 37.42518, 23.08245, 7.710317,
  -8.952087, -25.66975, -39.07905, -47.71579, -51.00347, -49.13211, -40.5117, 
    -26.77046, -13.02728, 0.05396039, 12.0524, 23.06087, 32.90032, 40.63223, 
    44.80841, 44.42027, 40.8101, 32.33792, 19.52864, 6.429458,
  -8.680319, -24.87808, -37.78508, -45.84899, -48.39751, -45.61121, 
    -37.03951, -24.15419, -10.58928, 2.929039, 15.67566, 27.23701, 36.93014, 
    43.4728, 45.28839, 41.5574, 34.15936, 25.06474, 14.7433, 4.757007,
  -8.367161, -23.98036, -36.36882, -43.89514, -45.73133, -41.92244, 
    -33.52592, -21.98254, -8.971597, 4.793093, 18.28484, 30.51069, 40.18296, 
    45.59449, 45.02596, 37.92479, 26.77305, 17.52895, 10.14617, 3.210453,
  -8.17645, -23.43475, -35.49448, -42.60479, -43.7156, -38.62022, -30.19488, 
    -20.06808, -7.788923, 5.942511, 19.85872, 32.45412, 41.90814, 46.19212, 
    43.61407, 34.04411, 20.42356, 11.81454, 7.147548, 2.280969,
  -8.222074, -23.5569, -35.60432, -42.45295, -42.83879, -36.36192, -27.44073, 
    -18.0592, -6.332018, 7.010953, 20.61958, 32.74601, 41.35553, 44.45808, 
    40.7781, 30.79415, 17.5272, 10.48608, 7.316301, 2.492983,
  -7.783059, -22.40804, -34.29367, -41.98576, -44.63146, -41.83231, 
    -35.57736, -24.53912, -6.84904, 14.84174, 37.58821, 58.18573, 73.28196, 
    79.76471, 75.53751, 60.69614, 38.38868, 19.36402, 8.88769, 2.456524,
  -8.353537, -24.05282, -36.81985, -45.13011, -48.23254, -46.15659, 
    -38.76635, -25.48749, -6.86278, 15.1569, 37.93541, 58.27677, 72.83444, 
    78.77555, 74.67533, 61.48814, 42.98889, 25.39217, 12.55283, 3.680161,
  -8.852053, -25.47714, -38.97097, -47.73624, -51.05746, -49.18595, 
    -41.14826, -26.75531, -7.553002, 14.83298, 37.89825, 58.44241, 73.09789, 
    79.0899, 75.17139, 62.56817, 45.37763, 28.11009, 14.12193, 4.189902,
  -7.564929, -21.65483, -32.76643, -39.46875, -41.16231, -38.06153, 
    -31.18344, -20.58916, -6.142004, 10.98142, 29.09966, 46.0606, 59.53432, 
    67.46596, 68.54298, 62.59012, 50.77349, 36.16738, 21.3623, 6.998292,
  -7.228909, -20.69444, -31.31371, -37.70515, -39.2724, -36.19323, -29.5204, 
    -19.28262, -5.265425, 11.34578, 28.88865, 45.26204, 58.23044, 65.8595, 
    66.92852, 61.25508, 49.85717, 35.71114, 21.25817, 6.99873,
  -6.89532, -19.71889, -29.77601, -35.73652, -37.03304, -33.8278, -27.33514, 
    -17.5553, -4.113688, 11.77329, 28.49198, 44.05666, 56.40401, 63.77009, 
    65.00415, 59.81119, 48.91588, 35.28028, 21.23863, 7.040614,
  -6.612323, -18.86744, -28.37156, -33.84493, -34.77104, -31.31235, 
    -24.96962, -15.71303, -2.92351, 12.10729, 27.82672, 42.42873, 54.09851, 
    61.28203, 62.86518, 58.32905, 47.9719, 34.82869, 21.22499, 7.090059,
  -6.364327, -18.09469, -27.03091, -31.95104, -32.41852, -28.62806, 
    -22.43289, -13.77041, -1.729493, 12.30029, 26.8377, 40.32782, 51.28363, 
    58.3895, 60.51345, 56.78559, 46.97291, 34.1973, 20.98363, 7.045365,
  -6.152084, -17.41649, -25.82574, -30.2443, -30.34912, -26.39354, -20.42057, 
    -12.33086, -1.0585, 11.9153, 25.19561, 37.56085, 47.9401, 55.28039, 
    58.35216, 55.75431, 46.55311, 33.77803, 20.55886, 6.876444,
  -7.002536, -19.74337, -29.02538, -33.47636, -32.68294, -27.04877, 
    -18.45868, -9.257074, -0.5703061, 7.536592, 14.84504, 21.29163, 26.88585, 
    31.50799, 34.74586, 35.97162, 35.10575, 30.97403, 21.66323, 7.707413,
  -7.738431, -21.89919, -32.52711, -38.36885, -39.1657, -35.35406, -26.75187, 
    -15.5193, -5.2751, 3.916564, 11.99589, 19.28349, 26.17193, 32.72108, 
    38.41271, 42.23374, 43.63003, 38.37428, 25.66404, 8.955738,
  -8.733225, -24.78973, -37.10385, -44.44256, -46.6473, -44.22988, -35.43698, 
    -22.33988, -10.43607, 0.2094415, 9.637213, 18.39761, 27.04028, 35.59348, 
    43.35806, 49.08753, 52.10927, 45.88302, 30.08752, 10.42105,
  -9.766819, -27.77761, -41.76472, -50.44027, -53.67297, -52.02555, 
    -42.88248, -28.27415, -14.75519, -2.454965, 8.662466, 19.1989, 29.67088, 
    39.94551, 49.11742, 55.79527, 59.33347, 52.0738, 33.87242, 11.69861,
  -10.57051, -30.06824, -45.22899, -54.6773, -58.29459, -56.73156, -47.13756, 
    -31.48958, -16.72513, -3.077574, 9.428221, 21.34755, 33.09036, 44.35406, 
    54.06894, 60.76306, 63.86197, 55.60496, 35.9774, 12.39417,
  -10.96969, -31.1578, -46.72089, -56.19806, -59.50245, -57.43431, -47.45782, 
    -31.43703, -16.06923, -1.691853, 11.58121, 24.19114, 36.40879, 47.79281, 
    57.16429, 63.01049, 64.83367, 55.70376, 35.82181, 12.29293,
  -10.99127, -31.14988, -46.47989, -55.44866, -58.00074, -55.09891, 
    -44.97556, -29.31502, -13.96331, 0.6672647, 14.33004, 27.24583, 39.46217, 
    50.3758, 58.7073, 62.91509, 62.59355, 52.64139, 33.58697, 11.46072,
  -10.79928, -30.54508, -45.36053, -53.64007, -55.30999, -51.42775, 
    -41.40977, -26.74988, -11.84061, 2.862056, 16.91883, 30.19571, 42.38081, 
    52.61573, 59.46698, 61.34868, 57.98034, 47.20903, 29.89803, 10.13695,
  -10.57625, -29.88047, -44.22331, -51.89633, -52.70943, -47.67823, -37.861, 
    -24.64393, -10.40161, 4.357369, 18.94847, 32.78287, 45.07676, 54.62046, 
    59.76488, 58.87062, 51.81361, 40.4199, 25.63107, 8.665152,
  -10.43863, -29.47854, -43.52624, -50.71486, -50.63114, -44.10755, 
    -34.34302, -22.77322, -9.2978, 5.441452, 20.49506, 34.81046, 47.11948, 
    55.855, 59.1887, 55.51762, 44.90794, 33.56332, 21.86731, 7.461738,
  -10.48378, -29.59258, -43.58868, -50.41114, -49.42835, -41.29688, 
    -31.25714, -20.8861, -7.951854, 6.655083, 21.77976, 36.05521, 47.89603, 
    55.55453, 57.26337, 51.73534, 39.29304, 29.18719, 20.36785, 7.162384,
  -10.14348, -28.80934, -43.02914, -51.0349, -52.23284, -46.75346, -38.63196, 
    -26.83722, -8.157217, 15.02581, 40.06341, 64.11121, 84.1581, 97.10458, 
    99.94078, 90.36871, 68.15321, 44.10655, 25.4877, 8.237379,
  -10.70087, -30.41879, -45.52647, -54.24634, -56.16267, -51.80383, 
    -42.81873, -28.67244, -8.628447, 15.42018, 41.04562, 65.34846, 85.19499, 
    97.55396, 99.92324, 91.04166, 71.9427, 49.41435, 28.78439, 9.371364,
  -11.23531, -31.92843, -47.77622, -56.97347, -59.22076, -55.33231, 
    -45.79887, -30.37882, -9.544452, 15.11085, 41.26616, 65.98538, 86.06307, 
    98.47115, 100.876, 92.38779, 74.59725, 52.41529, 30.46307, 9.913744,
  -8.494239, -24.20615, -36.35181, -43.41382, -44.92626, -41.30972, 
    -33.80649, -22.52917, -7.266226, 10.87612, 30.34416, 49.1347, 65.03026, 
    75.93987, 80.20532, 76.88354, 66.06374, 49.99686, 31.07979, 10.49668,
  -8.16336, -23.26265, -34.92728, -41.67978, -43.04647, -39.40307, -32.0317, 
    -21.0248, -6.108381, 11.58442, 30.50352, 48.68307, 63.98722, 74.43964, 
    78.49213, 75.24966, 64.72929, 49.12691, 30.68309, 10.39383,
  -7.85905, -22.36422, -33.48762, -39.79693, -40.84656, -36.9942, -29.67852, 
    -18.98084, -4.500469, 12.56923, 30.69829, 48.01707, 62.55446, 72.51817, 
    76.47762, 73.50397, 63.39552, 48.32286, 30.39865, 10.34316,
  -7.600342, -21.57788, -32.1705, -37.99306, -38.64757, -34.48728, -27.18815, 
    -16.82109, -2.809642, 13.55381, 30.76011, 47.08607, 60.79323, 70.31483, 
    74.3187, 71.75324, 62.09047, 47.50527, 30.08733, 10.28242,
  -7.346431, -20.79661, -30.84164, -36.15339, -36.39531, -31.93531, 
    -24.67432, -14.67371, -1.189859, 14.38301, 30.55866, 45.80859, 58.68278, 
    67.85754, 72.0548, 70.00581, 60.79575, 46.5443, 29.51843, 10.10489,
  -7.087369, -20.01376, -29.55719, -34.46979, -34.47702, -29.95576, 
    -22.84497, -13.19738, -0.2398546, 14.55419, 29.72175, 43.97574, 56.20686, 
    65.34088, 70.08508, 68.81374, 60.10277, 45.84526, 28.81256, 9.814613,
  -7.787515, -21.9286, -32.18693, -37.12155, -36.40686, -30.64425, -21.44046, 
    -10.86494, -0.5199575, 9.338877, 18.34647, 26.34244, 33.29684, 39.10695, 
    43.38816, 45.41963, 44.64835, 39.18663, 27.30172, 9.745531,
  -8.420586, -23.83658, -35.43184, -41.86179, -42.8544, -38.93263, -29.74736, 
    -17.21494, -5.254872, 5.856925, 15.83607, 24.80345, 33.03782, 40.60666, 
    47.0719, 51.40518, 52.5999, 46.05176, 31.00974, 10.88994,
  -9.28125, -26.37805, -39.56958, -47.53005, -50.03001, -47.60029, -38.29872, 
    -23.96217, -10.36374, 2.223083, 13.58104, 24.01242, 33.92733, 43.37651, 
    51.78076, 57.91409, 60.64509, 53.15667, 35.16147, 12.25602,
  -10.1683, -28.96715, -43.67755, -52.92695, -56.48821, -54.91537, -45.35638, 
    -29.62314, -14.56823, -0.496507, 12.39046, 24.45772, 36.10014, 47.23276, 
    57.08694, 64.28648, 67.69077, 59.26051, 38.88734, 13.51346,
  -10.8275, -30.85121, -46.54211, -56.45896, -60.38834, -58.96852, -49.08183, 
    -32.50719, -16.49076, -1.384317, 12.61034, 25.86403, 38.70681, 50.90802, 
    61.53136, 69.08394, 72.42641, 63.16255, 41.28213, 14.3206,
  -11.10261, -31.5796, -47.47233, -57.28279, -60.85202, -58.97966, -48.85722, 
    -32.16768, -15.90253, -0.4515765, 13.97614, 27.71235, 41.00316, 53.50465, 
    64.16311, 71.39543, 74.03667, 64.12557, 41.79358, 14.47211,
  -11.04203, -31.31808, -46.80238, -55.95832, -58.69905, -56.01414, 
    -45.87693, -29.8013, -13.90674, 1.397315, 15.85548, 29.66833, 42.93104, 
    55.18102, 65.27371, 71.55096, 72.80093, 62.33851, 40.52754, 14.00224,
  -10.82164, -30.60297, -45.44374, -53.76421, -55.51377, -51.82478, 
    -41.88105, -27.00388, -11.84529, 3.168897, 17.66599, 31.5849, 44.75013, 
    56.51306, 65.61483, 70.319, 69.36275, 58.34217, 37.90009, 13.0683,
  -10.61878, -29.96126, -44.25058, -51.82285, -52.57354, -47.66526, 
    -37.97285, -24.6825, -10.39337, 4.406911, 19.14986, 33.39792, 46.58803, 
    57.79443, 65.59084, 68.15157, 64.17411, 52.67743, 34.44044, 11.8874,
  -10.52895, -29.66148, -43.61253, -50.56391, -50.25116, -43.74612, 
    -34.16212, -22.66611, -9.257141, 5.396582, 20.47059, 35.10371, 48.29468, 
    58.79076, 64.97861, 64.9827, 57.52089, 46.00525, 30.83938, 10.74885,
  -10.62509, -29.89135, -43.76534, -50.23379, -48.86962, -40.65142, 
    -30.90888, -20.82848, -7.988945, 6.60154, 21.86705, 36.61343, 49.49873, 
    59.02515, 63.50352, 61.18627, 50.97146, 40.39445, 28.62238, 10.23102,
  -10.44169, -29.57192, -43.91986, -51.64062, -52.17226, -45.78354, 
    -37.31178, -25.89114, -7.670413, 15.25194, 40.44361, 65.27444, 86.97176, 
    102.6299, 109.1532, 103.4592, 83.55145, 58.85479, 36.32825, 12.2001,
  -11.04286, -31.31122, -46.63381, -55.16881, -56.53853, -51.3372, -42.1716, 
    -28.47085, -8.645677, 15.49434, 41.6636, 67.15557, 89.03288, 104.347, 
    110.3289, 104.7881, 87.05913, 63.45859, 39.19083, 13.19944,
  -11.60799, -32.90966, -49.02524, -58.09386, -59.87226, -55.23784, 
    -45.58967, -30.57445, -9.824021, 15.09699, 41.98839, 68.09582, 90.38704, 
    105.8709, 111.8908, 106.6071, 89.97675, 66.59045, 40.93722, 13.7667 ;

 hv =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -0.01967761, -0.4352752, -3.189604, -8.978535, -12.23629, 
    -12.74275, -12.76649, -12.76649, -12.76649, -12.76649, -12.76649, 
    -12.74275, -12.23629, -8.978535, -3.189604, -0.4352752, -0.01967761,
  0, 0, 0, -0.3526604, -4.027499, -20.60457, -53.77649, -74.18636, -78.80141, 
    -79.25483, -79.25483, -79.25483, -79.25483, -79.25483, -78.80141, 
    -74.18636, -53.77649, -20.60457, -4.027499, -0.3526604,
  0, 0, 0, -1.834447, -15.06886, -52.64848, -115.7051, -160.6247, -174.3762, 
    -176.0672, -176.0672, -176.0672, -176.0672, -176.0672, -174.3762, 
    -160.6247, -115.7051, -52.64848, -15.06886, -1.834447,
  0, 0, 0, -1.856916, -15.24033, -52.18017, -105.9627, -145.2902, -157.5199, 
    -159.1111, -159.1111, -159.1111, -159.1111, -159.1111, -157.5199, 
    -145.2902, -105.9627, -52.18017, -15.24033, -1.856916,
  0, 0, 0, -0.3764539, -4.343614, -21.30734, -39.22413, -55.17839, -60.08724, 
    -60.7706, -60.7706, -60.7706, -60.7706, -60.7706, -60.08724, -55.17839, 
    -39.22413, -21.30734, -4.343614, -0.3764539,
  0, 0, 0, -0.02100252, -0.4896586, -3.56352, -6.384347, -9.482255, 
    -10.46184, -10.58736, -10.58736, -10.58736, -10.58736, -10.58736, 
    -10.46184, -9.482255, -6.384347, -3.56352, -0.4896586, -0.02100252,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.02100252, 0.4896586, 3.56352, 6.384347, 9.482255, 10.46184, 
    10.58736, 10.58736, 10.58736, 10.58736, 10.58736, 10.46184, 9.482255, 
    6.384347, 3.56352, 0.4896586, 0.02100252,
  0, 0, 0, 0.3764539, 4.343614, 21.30734, 39.22413, 55.17839, 60.08724, 
    60.7706, 60.7706, 60.7706, 60.7706, 60.7706, 60.08724, 55.17839, 
    39.22413, 21.30734, 4.343614, 0.3764539,
  0, 0, 0, 1.856916, 15.24033, 52.18017, 105.9627, 145.2902, 157.5199, 
    159.1111, 159.1111, 159.1111, 159.1111, 159.1111, 157.5199, 145.2902, 
    105.9627, 52.18017, 15.24033, 1.856916,
  0, 0, 0, 1.834447, 15.06886, 52.64848, 115.7051, 160.6247, 174.3762, 
    176.0672, 176.0672, 176.0672, 176.0672, 176.0672, 174.3762, 160.6247, 
    115.7051, 52.64848, 15.06886, 1.834447,
  0, 0, 0, 0.3526604, 4.027499, 20.60457, 53.77649, 74.18636, 78.80141, 
    79.25483, 79.25483, 79.25483, 79.25483, 79.25483, 78.80141, 74.18636, 
    53.77649, 20.60457, 4.027499, 0.3526604,
  0, 0, 0, 0.01967761, 0.4352752, 3.189604, 8.978535, 12.23629, 12.74275, 
    12.76649, 12.76649, 12.76649, 12.76649, 12.76649, 12.74275, 12.23629, 
    8.978535, 3.189604, 0.4352752, 0.01967761,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -1.483982e-05, -0.0006924636, -0.01148862, -0.0959114, -0.4257405, 
    -1.000566, -1.37499, -1.4755, -1.488466, -1.489292, -1.489306, -1.489292, 
    -1.488466, -1.4755, -1.37499, -1.000566, -0.4257405, -0.09594109, 
    -0.01216626,
  0, -0.0006084327, -0.01724106, -0.1923154, -1.162245, -4.401885, -10.06473, 
    -13.97968, -15.22131, -15.44909, -15.4706, -15.47138, -15.4706, 
    -15.44909, -15.22131, -13.97968, -10.06473, -4.401885, -1.162862, 
    -0.2095801,
  0, -0.008703556, -0.1650957, -1.322362, -6.125233, -19.32378, -41.89001, 
    -58.61727, -64.95157, -66.49261, -66.70441, -66.71632, -66.70441, 
    -66.49261, -64.95157, -58.61727, -41.89001, -19.32378, -6.134124, 
    -1.488657,
  0, -0.05843922, -0.8130453, -5.048312, -18.58049, -47.14565, -92.03905, 
    -128.6163, -144.9926, -149.9001, -150.7979, -150.8723, -150.7979, 
    -149.9001, -144.9926, -128.6163, -92.03905, -47.14565, -18.64234, 
    -5.879325,
  0, -0.1788347, -2.24571, -12.11221, -36.54682, -72.90214, -121.4297, 
    -171.7994, -197.6343, -205.9349, -207.51, -207.6383, -207.51, -205.9349, 
    -197.6343, -171.7994, -121.4297, -72.90214, -36.74054, -14.4527,
  0, -0.1815949, -2.307876, -12.45412, -36.92601, -72.47871, -110.6728, 
    -155.424, -177.9213, -185.3119, -186.7773, -186.9032, -186.7773, 
    -185.3119, -177.9213, -155.424, -110.6728, -72.47871, -37.1244, -14.88314,
  0, -0.06181528, -0.8968709, -5.607738, -19.71992, -47.10022, -65.76106, 
    -91.9437, -104.8842, -109.4054, -110.3811, -110.474, -110.3811, 
    -109.4054, -104.8842, -91.9437, -65.76106, -47.10022, -19.79486, -6.583194,
  0, -0.009371349, -0.1881541, -1.537523, -6.814981, -19.85835, -26.54994, 
    -38.21181, -44.16817, -46.25867, -46.70958, -46.75299, -46.70958, 
    -46.25867, -44.16817, -38.21181, -26.54994, -19.85835, -6.829762, 
    -1.750755,
  0, -0.0006677921, -0.01976805, -0.2308211, -1.364896, -4.768666, -6.146877, 
    -9.226855, -10.89776, -11.47999, -11.60295, -11.61462, -11.60295, 
    -11.47999, -10.89776, -9.226855, -6.146877, -4.768681, -1.366762, 
    -0.2544015,
  0, -2.225974e-05, -0.0007812203, -0.01395897, -0.1209926, -0.4899727, 
    -0.600044, -0.9434834, -1.145593, -1.216492, -1.231321, -1.232733, 
    -1.231321, -1.216492, -1.145593, -0.9434834, -0.600044, -0.4899876, 
    -0.1211316, -0.01495462,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 2.225974e-05, 0.0007812203, 0.01395897, 0.1209926, 0.4899727, 0.600044, 
    0.9434834, 1.145593, 1.216492, 1.231321, 1.232733, 1.231321, 1.216492, 
    1.145593, 0.9434834, 0.600044, 0.4899876, 0.1211316, 0.01495462,
  0, 0.0006677921, 0.01976805, 0.2308211, 1.364896, 4.768666, 6.146877, 
    9.226855, 10.89776, 11.47999, 11.60295, 11.61462, 11.60295, 11.47999, 
    10.89776, 9.226855, 6.146877, 4.768681, 1.366762, 0.2544015,
  0, 0.009371349, 0.1881541, 1.537523, 6.814981, 19.85835, 26.54994, 
    38.21181, 44.16817, 46.25867, 46.70958, 46.75299, 46.70958, 46.25867, 
    44.16817, 38.21181, 26.54994, 19.85835, 6.829762, 1.750755,
  0, 0.06181528, 0.8968709, 5.607738, 19.71992, 47.10022, 65.76106, 91.9437, 
    104.8842, 109.4054, 110.3811, 110.474, 110.3811, 109.4054, 104.8842, 
    91.9437, 65.76106, 47.10022, 19.79486, 6.583194,
  0, 0.1815949, 2.307876, 12.45412, 36.92601, 72.47871, 110.6728, 155.424, 
    177.9213, 185.312, 186.7773, 186.9032, 186.7773, 185.312, 177.9213, 
    155.424, 110.6728, 72.47871, 37.1244, 14.88314,
  0, 0.1788347, 2.24571, 12.11221, 36.54682, 72.90214, 121.4297, 171.7994, 
    197.6343, 205.9349, 207.51, 207.6383, 207.51, 205.9349, 197.6343, 
    171.7994, 121.4297, 72.90214, 36.74054, 14.4527,
  0, 0.05843922, 0.8128598, 5.04214, 18.50693, 46.74843, 91.0472, 127.273, 
    143.5746, 148.4756, 149.3733, 149.4477, 149.3733, 148.4756, 143.5746, 
    127.273, 91.0472, 46.74843, 18.56879, 5.872967,
  0, 0.008718396, 0.1598247, 1.211825, 5.22438, 15.20167, 31.64315, 44.40736, 
    49.71704, 51.11913, 51.32398, 51.3359, 51.32398, 51.11913, 49.71704, 
    44.40736, 31.64315, 15.20167, 5.233301, 1.372844,
  -3.115998e-05, -0.0006349122, -0.007029435, -0.04804701, -0.2179819, 
    -0.6740727, -1.379691, -1.905609, -2.114703, -2.166541, -2.174676, 
    -2.175414, -2.174676, -2.166541, -2.114703, -1.905609, -1.379691, 
    -0.6740991, -0.2186203, -0.05509306,
  -0.0005872581, -0.008844592, -0.07591648, -0.4220298, -1.634155, -4.621918, 
    -9.284207, -12.91608, -14.50535, -14.97279, -15.06438, -15.0749, 
    -15.06438, -14.97279, -14.50535, -12.91608, -9.284222, -4.622535, 
    -1.643124, -0.4982549,
  -0.005982158, -0.06722611, -0.4605001, -2.09819, -6.850674, -17.15917, 
    -33.10582, -46.26136, -52.73093, -55.00878, -55.56522, -55.64564, 
    -55.56522, -55.00878, -52.73093, -46.26136, -33.10606, -17.16538, 
    -6.920571, -2.565397,
  -0.03577322, -0.3210921, -1.810211, -6.878673, -18.93729, -40.85399, 
    -73.31889, -101.9884, -117.7118, -124.1855, -126.1142, -126.4546, 
    -126.1142, -124.1855, -117.7118, -101.9884, -73.3208, -40.89229, 
    -19.28307, -8.751168,
  -0.1341243, -1.017745, -4.904755, -15.88542, -36.90208, -66.92298, 
    -107.685, -149.2033, -174.322, -185.8486, -189.8159, -190.6237, 
    -189.8159, -185.8486, -174.322, -149.2033, -107.6931, -67.06528, 
    -38.02411, -21.077,
  -0.2993702, -2.134641, -9.483485, -27.30637, -54.24198, -82.73222, 
    -115.6348, -164.2644, -196.2919, -211.2443, -216.364, -217.3799, 
    -216.364, -211.2443, -196.2919, -164.2644, -115.6481, -83.02856, 
    -56.58631, -37.50962,
  -0.3068463, -2.214623, -9.870452, -28.08919, -54.78616, -83.333, -107.013, 
    -152.3438, -181.0006, -194.3422, -199.0037, -199.9547, -199.0037, 
    -194.3422, -181.0006, -152.3438, -107.0229, -83.6244, -57.20464, -38.78065,
  -0.1450774, -1.142517, -5.571281, -17.49569, -38.3326, -66.91639, 
    -79.95293, -111.3102, -130.3427, -139.6479, -143.159, -143.9356, 
    -143.159, -139.6479, -130.3427, -111.3102, -79.95815, -67.07035, 
    -39.67638, -23.76137,
  -0.03995442, -0.3771228, -2.167192, -7.945868, -20.13055, -40.12679, 
    -45.63746, -64.02128, -75.48746, -81.22345, -83.42668, -83.92268, 
    -83.42668, -81.22345, -75.48746, -64.02128, -45.64022, -40.18703, 
    -20.65032, -10.51619,
  -0.006784982, -0.08092504, -0.5714331, -2.533243, -7.57017, -17.05777, 
    -18.69564, -26.85381, -32.22659, -34.94556, -35.98455, -36.21709, 
    -35.98455, -34.94556, -32.22659, -26.85381, -18.69691, -17.07789, 
    -7.715024, -3.252907,
  -0.0006798548, -0.01072763, -0.09635334, -0.5305488, -1.8966, -4.741883, 
    -4.986995, -7.393084, -9.09621, -9.971436, -10.30355, -10.3771, 
    -10.30355, -9.971436, -9.09621, -7.393084, -4.987442, -4.747379, 
    -1.925232, -0.66006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0006798548, 0.01072763, 0.09635334, 0.5305488, 1.8966, 4.741883, 
    4.986995, 7.393084, 9.09621, 9.971436, 10.30355, 10.3771, 10.30355, 
    9.971436, 9.09621, 7.393084, 4.987442, 4.747379, 1.925232, 0.66006,
  0.006784982, 0.08092504, 0.5714331, 2.533243, 7.57017, 17.05777, 18.69564, 
    26.85381, 32.22659, 34.94556, 35.98455, 36.21709, 35.98455, 34.94556, 
    32.22659, 26.85381, 18.69691, 17.07789, 7.715024, 3.252907,
  0.03995442, 0.3771228, 2.167192, 7.945868, 20.13055, 40.12679, 45.63746, 
    64.02128, 75.48746, 81.22345, 83.42668, 83.92268, 83.42668, 81.22345, 
    75.48746, 64.02128, 45.64022, 40.18703, 20.65032, 10.51619,
  0.1450774, 1.142517, 5.571281, 17.49569, 38.3326, 66.91639, 79.95293, 
    111.3102, 130.3427, 139.6479, 143.159, 143.9356, 143.159, 139.6479, 
    130.3427, 111.3102, 79.95815, 67.07035, 39.67638, 23.76137,
  0.3068463, 2.214623, 9.870287, 28.08728, 54.77382, 83.28805, 106.937, 
    152.2483, 180.8996, 194.2395, 198.9001, 199.8509, 198.9001, 194.2395, 
    180.8996, 152.2483, 106.947, 83.57942, 57.19228, 38.77858,
  0.2993702, 2.134387, 9.479324, 27.26966, 54.04502, 82.06366, 114.2648, 
    162.447, 194.3237, 209.2422, 214.3558, 215.3709, 214.3558, 209.2422, 
    194.3237, 162.447, 114.2781, 82.35997, 56.38905, 37.46868,
  0.1340187, 1.014081, 4.859879, 15.5732, 35.50092, 62.56506, 98.64243, 
    136.804, 160.6281, 171.8253, 175.7398, 176.543, 175.7398, 171.8253, 
    160.6281, 136.804, 98.65056, 62.70728, 36.61928, 20.71971,
  0.03467194, 0.2934625, 1.537584, 5.325634, 13.05811, 24.53671, 39.96621, 
    55.15968, 64.97887, 69.67726, 71.2592, 71.5628, 71.2592, 69.67726, 
    64.97887, 55.15968, 39.96812, 24.57379, 13.37474, 6.920507,
  -0.01966096, -0.09356984, -0.3769259, -1.179819, -2.947691, -6.071634, 
    -10.38537, -14.29962, -16.74257, -17.90333, -18.32076, -18.41248, 
    -18.32076, -17.90335, -16.74258, -14.29987, -10.38795, -6.090291, 
    -3.04485, -1.563468,
  -0.1091148, -0.45707, -1.667758, -4.798502, -11.18117, -21.9226, -36.8447, 
    -50.70459, -59.63452, -64.16044, -65.93974, -66.36417, -65.93974, 
    -64.16045, -59.63464, -50.70643, -36.86172, -22.02942, -11.6717, -6.527561,
  -0.4162928, -1.499078, -4.801309, -12.19682, -25.24188, -44.65398, 
    -70.91399, -96.61977, -114.2228, -124.0557, -128.4238, -129.5773, 
    -128.4238, -124.0557, -114.2235, -96.6291, -70.989, -45.06735, -26.90721, 
    -17.30886,
  -1.202267, -3.771812, -10.65109, -23.80614, -43.25719, -67.73132, 
    -99.34253, -133.9255, -158.9665, -174.0664, -181.4854, -183.6113, 
    -181.4854, -174.0665, -158.9692, -133.957, -99.57255, -68.89642, 
    -47.51942, -35.43961,
  -2.655507, -7.442234, -18.79523, -37.2428, -59.60435, -82.55583, -109.7858, 
    -148.8952, -178.8301, -197.5724, -207.2679, -210.168, -207.2679, 
    -197.5727, -178.836, -148.9632, -110.2753, -84.98074, -67.94872, -58.1062,
  -4.413054, -11.66492, -27.3123, -49.15438, -70.62638, -88.07574, -103.6437, 
    -146.2946, -181.0816, -202.7178, -213.5979, -216.7706, -213.5979, 
    -202.7178, -181.0847, -146.357, -104.2939, -91.82533, -83.40381, -79.66093,
  -4.627999, -12.25616, -28.40728, -50.35893, -71.88005, -90.65296, 
    -98.16039, -140.644, -173.6034, -193.6101, -203.6196, -206.5501, 
    -203.6196, -193.6101, -173.6045, -140.6816, -98.6809, -94.43188, 
    -85.12518, -82.11523,
  -3.053598, -8.605544, -21.11578, -39.88051, -61.61316, -85.45752, 
    -88.11773, -122.3865, -146.9796, -162.1615, -170.1346, -172.5728, 
    -170.1346, -162.1616, -146.9813, -122.4149, -88.43169, -88.07407, 
    -71.2997, -64.14575,
  -1.4704, -4.64545, -12.58385, -26.06817, -44.04706, -66.62708, -65.66868, 
    -89.9291, -107.3878, -118.4709, -124.4421, -126.2993, -124.4421, 
    -118.471, -107.3895, -89.95163, -65.8717, -68.12051, -49.7962, -41.23493,
  -0.5302659, -1.931299, -5.911335, -13.66947, -25.39493, -41.46014, 
    -39.53369, -54.15867, -65.08859, -72.18568, -76.04588, -77.25049, 
    -76.04588, -72.18573, -65.08995, -54.17506, -39.65553, -42.19461, 
    -28.1728, -21.25537,
  -0.1393122, -0.5896105, -2.046163, -5.276791, -10.69323, -18.53415, 
    -17.24325, -23.82448, -28.97532, -32.37799, -34.23338, -34.81137, 
    -34.23338, -32.37801, -28.97605, -23.83302, -17.29958, -18.82054, 
    -11.70849, -8.075982,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.1393122, 0.5896105, 2.046163, 5.276791, 10.69323, 18.53415, 17.24325, 
    23.82448, 28.97532, 32.37799, 34.23338, 34.81137, 34.23338, 32.37801, 
    28.97605, 23.83302, 17.29958, 18.82054, 11.70849, 8.075982,
  0.5302659, 1.931299, 5.911328, 13.66931, 25.3943, 41.45872, 39.53278, 
    54.15767, 65.08747, 72.18443, 76.04454, 77.24911, 76.04454, 72.18447, 
    65.08884, 54.17405, 39.65461, 42.19315, 28.17214, 21.25517,
  1.470397, 4.645368, 12.58316, 26.06443, 44.03379, 66.59633, 65.6452, 
    89.90311, 107.36, 118.441, 124.4104, 126.2668, 124.4104, 118.441, 
    107.3617, 89.92564, 65.84805, 68.08932, 49.78239, 41.23018,
  3.053459, 8.604194, 21.10696, 39.84033, 61.48149, 85.1454, 87.80979, 
    122.0335, 146.6104, 161.7764, 169.7356, 172.1684, 169.7356, 161.7764, 
    146.6121, 122.0616, 88.1224, 87.75959, 71.16455, 64.09543,
  4.626396, 12.2443, 28.34113, 50.09068, 71.06482, 88.75107, 95.37286, 
    137.1197, 169.759, 189.6266, 199.5699, 202.4792, 199.5699, 189.6266, 
    169.7599, 137.1565, 95.89089, 92.5254, 84.29547, 81.77927,
  4.40161, 11.59417, 26.96925, 47.91492, 67.18579, 80.49397, 90.69651, 
    129.0716, 161.5332, 182.1638, 192.6968, 195.7924, 192.6968, 182.1638, 
    161.5363, 129.1338, 91.34564, 84.23224, 79.88959, 78.07276,
  2.598127, 7.139299, 17.5099, 33.11758, 49.2465, 61.31767, 73.65694, 
    99.73178, 121.8525, 136.9206, 145.2861, 147.8915, 145.2861, 136.9209, 
    121.8584, 99.79991, 74.14144, 63.68769, 57.26694, 52.64904,
  0.994446, 2.807955, 7.030467, 13.49411, 20.14011, 24.64341, 28.69061, 
    36.62458, 44.51564, 50.88948, 54.86453, 56.17401, 54.86453, 50.8896, 
    44.51835, 36.65439, 28.89244, 25.58883, 23.30685, 21.23963,
  -0.4314921, -1.053732, -2.585984, -5.401428, -9.676617, -15.37907, 
    -22.53586, -29.93905, -35.95074, -40.04436, -42.27036, -42.95354, 
    -42.27042, -40.04488, -35.95486, -29.96367, -22.64785, -15.78021, 
    -10.83754, -8.17095,
  -1.555897, -3.560417, -8.291697, -16.57647, -28.59911, -44.16745, -63.9051, 
    -84.66095, -101.2172, -112.474, -118.6975, -120.6419, -118.6978, 
    -112.4765, -101.2353, -84.76136, -64.33485, -45.62964, -32.6222, -25.67388,
  -3.841238, -7.878544, -16.58271, -30.14957, -47.54357, -67.84286, 
    -93.02544, -121.6876, -144.9855, -161.3947, -170.94, -174.039, -170.9408, 
    -161.4025, -145.0389, -121.9619, -94.12209, -71.342, -56.49863, -48.74403,
  -7.744346, -14.2461, -26.91326, -44.10515, -62.98735, -82.28612, -105.278, 
    -137.3047, -164.0572, -183.3577, -194.9856, -198.8604, -194.9876, 
    -183.3753, -164.1718, -137.8719, -107.4555, -88.92289, -78.90563, 
    -74.62518,
  -13.01255, -21.80302, -37.34991, -55.73774, -72.88318, -87.98985, 
    -103.3885, -137.3527, -166.8448, -188.2277, -201.1682, -205.4982, 
    -201.1709, -188.2526, -167.0135, -138.2253, -106.8309, -98.3769, 
    -96.52946, -98.2122,
  -18.3113, -28.93774, -46.24686, -64.29873, -78.51865, -89.06976, -93.45741, 
    -129.9515, -163.688, -188.2654, -202.8774, -207.6952, -202.8776, 
    -188.2716, -163.7772, -130.7362, -97.65998, -102.882, -109.1364, -117.0216,
  -19.38282, -30.29923, -47.77475, -65.90646, -80.75799, -93.02949, -89.6151, 
    -127.377, -160.942, -184.653, -198.4808, -203.0054, -198.4802, -184.6518, 
    -160.9755, -127.9028, -93.23457, -107.2222, -112.4886, -120.3423,
  -15.33649, -24.85142, -40.78598, -58.9807, -76.68929, -94.74299, -88.1214, 
    -121.9271, -149.1373, -167.9014, -178.932, -182.5856, -178.9325, 
    -167.9064, -149.1834, -122.3117, -90.5778, -106.15, -103.2833, -106.0895,
  -9.862552, -17.17246, -30.15956, -46.36507, -64.0498, -84.18932, -75.72521, 
    -102.3277, -122.9761, -137.357, -145.9618, -148.8442, -145.9625, 
    -137.3635, -123.0236, -102.6381, -77.46306, -92.13487, -83.45133, 
    -82.22791,
  -5.154963, -9.836667, -18.72212, -30.72789, -44.87181, -61.95649, 
    -54.45384, -72.46506, -86.48517, -96.42078, -102.4442, -104.4748, 
    -102.4448, -96.42688, -86.52757, -72.70743, -55.60136, -66.7651, 
    -56.96598, -53.96564,
  -2.022524, -4.21454, -8.621619, -14.94755, -22.75967, -32.47306, -28.17188, 
    -37.23159, -44.38913, -49.52673, -52.6623, -53.7221, -52.66272, 
    -49.53051, -44.41462, -37.36828, -28.74902, -34.69686, -28.41808, 
    -26.11248,
  0, -1.832988e-05, -9.19906e-05, -0.0002882203, -0.0007579019, -0.001270073, 
    -0.0006334081, -0.0006388605, -0.0007077602, -0.0008190513, -0.000928168, 
    -0.0009409337, -0.0009262228, -0.0008504329, -0.0007314094, 
    -0.0006360859, -0.0006712821, -0.001366725, -0.0008976159, -0.0004774202,
  2.022485, 4.214312, 8.620529, 14.94376, 22.75022, 32.45689, 28.16303, 
    37.22255, 44.37935, 49.51585, 52.65041, 53.7098, 52.65085, 49.51962, 
    44.40481, 37.35911, 28.73972, 34.6796, 28.4073, 26.10678,
  5.15448, 9.83431, 18.71235, 30.69703, 44.79758, 61.82483, 54.37125, 
    72.37904, 86.39494, 96.32354, 102.3401, 104.3679, 102.3408, 96.32964, 
    86.43713, 72.62025, 55.51524, 66.62663, 56.88352, 53.9209,
  9.858662, 17.15587, 30.09779, 46.18456, 63.63047, 83.41595, 75.14016, 
    101.692, 122.3197, 136.6687, 145.2406, 148.1093, 145.2413, 136.675, 
    122.3659, 101.9958, 76.86031, 91.33581, 82.99715, 81.97394,
  15.31351, 24.76542, 40.49386, 58.18314, 74.90208, 91.38754, 84.87765, 
    118.1409, 145.1564, 163.7849, 174.7006, 178.3071, 174.701, 163.789, 
    145.1971, 118.5034, 87.28777, 102.7351, 101.3809, 104.9824,
  19.27924, 29.95493, 46.70147, 63.16828, 74.91741, 82.32845, 75.40214, 
    109.3603, 140.6933, 163.1974, 176.4305, 180.774, 176.4296, 163.194, 
    140.7166, 109.8595, 78.98038, 96.41237, 106.2853, 116.5115,
  17.94107, 27.83792, 43.11051, 56.90223, 63.84209, 63.75068, 55.7999, 
    80.59065, 105.9238, 125.4296, 137.5536, 141.652, 137.5536, 125.4356, 
    106.0133, 81.37375, 59.94393, 77.23277, 93.27911, 106.3315,
  11.95066, 18.98075, 30.03004, 39.92233, 44.02488, 41.72474, 35.79807, 
    48.07859, 61.07509, 71.87806, 79.30221, 81.97462, 79.30506, 71.90365, 
    61.24364, 48.92374, 39.02197, 51.12419, 64.49316, 74.40536,
  5.275858, 8.328547, 12.98213, 16.73679, 17.55274, 15.41305, 11.98952, 
    13.42739, 16.05498, 19.26197, 22.09078, 23.23384, 22.09291, 19.27935, 
    16.15731, 13.88429, 13.56603, 19.69898, 26.56513, 31.45946,
  -1.616347, -2.927933, -5.623295, -9.619379, -14.53404, -20.01976, 
    -26.44032, -33.60443, -40.14002, -45.36613, -48.72733, -49.88239, 
    -48.72858, -45.37429, -40.181, -33.76944, -26.98001, -21.47935, 
    -17.83056, -15.89524,
  -4.995333, -8.682455, -16.08485, -26.75149, -39.54997, -53.75935, 
    -70.91273, -90.71545, -108.0423, -121.3633, -129.7372, -132.588, 
    -129.7418, -121.3913, -108.1779, -91.24451, -72.60015, -58.22865, 
    -49.41294, -45.01262,
  -10.29419, -16.3656, -27.74697, -42.7051, -59.01087, -75.87485, -96.02972, 
    -122.2174, -145.0799, -162.6191, -173.7447, -177.5656, -173.756, 
    -162.685, -145.3827, -123.3479, -99.47464, -84.59035, -77.22028, -74.38605,
  -17.68888, -25.61255, -39.34595, -55.54596, -71.23993, -86.0849, -102.818, 
    -131.5975, -157.0064, -176.421, -188.7776, -193.0397, -188.798, 
    -176.5373, -157.5316, -133.5267, -108.5462, -100.0256, -98.7162, -100.3391,
  -26.24641, -35.06928, -49.34585, -64.59894, -77.6826, -88.85964, -98.15033, 
    -128.7441, -156.6374, -177.906, -191.3559, -195.9768, -191.3792, 
    -178.0452, -157.3061, -131.3568, -106.197, -108.2024, -113.9242, -120.5283,
  -34.15342, -43.28815, -57.28482, -70.96098, -81.2177, -88.90116, -87.99879, 
    -120.8196, -152.7528, -177.6125, -193.2884, -198.6387, -193.2891, 
    -177.6486, -153.129, -123.2147, -97.52266, -113.0303, -124.9908, -136.0393,
  -36.11758, -45.1267, -58.99994, -72.86086, -83.94222, -93.24969, -84.58889, 
    -118.871, -151.3572, -175.9643, -191.1251, -196.2386, -191.1196, 
    -175.9577, -151.5228, -120.6162, -93.13844, -118.2218, -129.2316, 
    -139.8528,
  -30.82481, -39.35496, -53.14719, -68.32803, -82.69075, -97.23336, 
    -85.58342, -117.6883, -145.1824, -165.0318, -177.0464, -181.0848, 
    -177.0494, -165.0556, -145.3672, -118.9648, -91.79398, -118.5693, 
    -122.6621, -129.0041,
  -22.4169, -29.9819, -42.65755, -57.50555, -72.93433, -90.12621, -77.36586, 
    -103.8758, -125.2004, -140.3824, -149.6082, -152.7252, -149.6134, 
    -140.4147, -125.3826, -104.8715, -81.93837, -106.2207, -104.3755, 
    -106.9457,
  -13.65554, -19.37174, -29.21103, -41.20493, -54.31033, -69.64004, 
    -58.84336, -77.43696, -91.99219, -102.3887, -108.7634, -110.929, 
    -108.7687, -102.4205, -92.1549, -78.19437, -61.92916, -80.1694, 
    -75.62405, -75.86172,
  -6.199827, -9.27584, -14.66981, -21.40092, -28.9359, -37.94138, -31.79585, 
    -41.33949, -48.75843, -54.08823, -57.37619, -58.49675, -57.37957, 
    -54.10825, -48.85698, -41.76331, -33.36911, -43.10594, -39.62846, 
    -39.20385,
  -0.0001616009, -0.0006870263, -0.002413273, -0.006616501, -0.01394199, 
    -0.02097762, -0.01044726, -0.01010023, -0.01075009, -0.01190138, 
    -0.01300092, -0.01344548, -0.01300261, -0.01195235, -0.01087956, 
    -0.01050257, -0.01162673, -0.02357849, -0.01714141, -0.01101734,
  6.198302, 9.270499, 14.65267, 21.35667, 28.84531, 37.80112, 31.7185, 
    41.26303, 48.67928, 54.0033, 57.28533, 58.40341, 57.28871, 54.02316, 
    48.77704, 41.68382, 33.2842, 42.95171, 39.52097, 39.13393,
  13.64575, 19.34138, 29.12113, 40.98582, 53.87171, 68.93262, 58.39304, 
    76.97344, 91.52118, 101.8972, 108.2486, 110.404, 108.2538, 101.9283, 
    91.6797, 77.71496, 61.44427, 79.41161, 75.12131, 75.53012,
  22.36822, 29.84497, 42.27996, 56.62936, 71.21294, 87.24677, 75.15421, 
    101.4478, 122.7172, 137.834, 146.985, 150.0686, 146.9896, 137.8626, 
    122.8815, 102.3843, 79.6185, 103.2101, 102.4537, 105.6538,
  30.63168, 38.858, 51.86532, 65.49608, 77.27531, 88.07832, 76.7588, 
    107.1919, 133.9679, 153.4331, 165.1955, 169.1381, 165.1963, 153.4452, 
    134.1051, 108.3449, 82.78749, 109.1559, 116.6858, 124.8481,
  35.49193, 43.6497, 55.43985, 65.42706, 70.37055, 71.03877, 56.71862, 
    83.70975, 111.1941, 132.7325, 146.2817, 150.8959, 146.2719, 132.7071, 
    111.3052, 85.35684, 65.11466, 95.46724, 114.1199, 128.7402,
  32.4608, 39.63277, 49.1257, 55.09956, 54.22577, 47.4825, 31.23871, 
    47.92695, 66.71502, 82.3781, 92.83972, 96.52863, 92.8401, 82.41534, 
    67.0974, 50.28329, 40.37428, 70.13341, 93.98781, 111.3467,
  22.4197, 27.53863, 33.91246, 36.92064, 34.20124, 26.81624, 14.88528, 
    21.57127, 29.29796, 35.88723, 40.6101, 42.36097, 40.63455, 36.02817, 
    29.94437, 23.97056, 21.89285, 42.74533, 61.88435, 75.46671,
  10.3883, 12.50472, 14.80353, 15.18251, 13.02199, 9.193375, 4.214333, 
    3.842202, 4.148524, 4.908947, 5.824281, 6.241668, 5.845121, 5.014826, 
    4.572361, 5.217303, 7.797578, 16.71661, 25.45004, 31.5456,
  -4.155516, -6.001171, -9.320594, -13.40651, -17.46109, -21.13637, 
    -25.11554, -30.12932, -35.09414, -39.52146, -42.68213, -43.84025, 
    -42.69437, -39.57714, -35.2982, -30.75492, -26.73075, -24.68821, 
    -24.11867, -24.06852,
  -11.64892, -16.40551, -24.89182, -35.28617, -45.68726, -55.51822, 
    -66.93584, -82.29556, -96.58566, -108.4365, -116.4638, -119.3279, 
    -116.4987, -108.5927, -97.15352, -84.0294, -71.3875, -65.26128, 
    -63.79477, -63.95656,
  -21.14554, -27.79282, -39.17209, -52.39684, -65.01498, -76.7477, -90.29829, 
    -111.9302, -131.704, -147.6015, -158.1467, -161.8744, -158.2155, 
    -147.9002, -132.7625, -115.0809, -98.13513, -93.29594, -94.4325, -96.91576,
  -32.25516, -39.3486, -51.00818, -63.85151, -75.43525, -85.92162, -96.63938, 
    -121.6599, -144.5016, -162.4554, -174.173, -178.2867, -174.2762, 
    -162.9029, -146.0878, -126.3669, -108.1528, -109.4122, -115.0757, 
    -120.8406,
  -43.54517, -49.87896, -60.10515, -70.99532, -80.26163, -88.31161, 
    -92.48969, -119.8458, -145.5252, -165.6944, -178.7688, -183.3347, 
    -178.8714, -166.1724, -147.3593, -125.6953, -107.3792, -118.2641, 
    -128.5189, -137.3906,
  -53.31684, -58.57009, -67.08752, -75.90469, -82.77866, -88.30913, 
    -83.24112, -112.7426, -142.3126, -166.3591, -182.1003, -187.5802, 
    -182.1034, -166.4996, -143.4411, -118.2584, -100.475, -124.0105, 
    -138.4145, -150.0762,
  -56.09715, -60.82433, -68.95916, -77.95675, -85.62127, -92.51997, 
    -79.93871, -110.758, -141.2242, -165.5154, -181.0495, -186.3783, 
    -181.0234, -165.5064, -141.8155, -115.0932, -95.88755, -129.553, 
    -143.0037, -154.0514,
  -50.3123, -55.19492, -64.11944, -74.9504, -85.69741, -96.91197, -81.46574, 
    -111.0079, -137.5991, -157.5285, -169.8096, -173.9623, -169.8178, 
    -157.6001, -138.1463, -114.2328, -93.68, -129.7687, -137.8416, -145.5426,
  -39.70232, -44.69962, -53.87405, -65.31322, -77.45388, -91.11656, 
    -75.20201, -100.4082, -121.3526, -136.4348, -145.5949, -148.6842, 
    -145.6134, -136.5298, -121.838, -102.8362, -84.46918, -117.1122, 
    -120.1378, -124.731,
  -26.67191, -30.98928, -38.80568, -48.56029, -59.20398, -71.65968, 
    -58.56627, -76.65089, -90.88311, -100.9503, -107.0594, -109.1252, 
    -107.0794, -101.045, -91.2952, -78.4015, -64.88788, -89.42168, -89.30528, 
    -91.57887,
  -13.195, -15.74369, -20.29732, -25.94997, -32.17586, -39.58517, -32.18391, 
    -41.5499, -48.72246, -53.76814, -56.83757, -57.87838, -56.85044, 
    -53.82799, -48.96806, -42.50053, -35.41702, -48.56715, -47.7244, -48.57841,
  -0.00353562, -0.009418536, -0.02474869, -0.05448993, -0.09842989, 
    -0.1380206, -0.06995916, -0.06583223, -0.06679557, -0.0706763, 
    -0.07494253, -0.0767677, -0.07501744, -0.07112705, -0.06858969, 
    -0.07162303, -0.08223195, -0.1601351, -0.125245, -0.09268969,
  13.17511, 15.69523, 20.17747, 25.696, 31.72315, 38.92987, 31.81577, 
    41.19084, 48.36434, 53.39886, 56.45338, 57.48744, 56.46584, 53.45644, 
    48.60054, 42.11276, 34.99466, 47.82976, 47.16976, 48.16631,
  26.58704, 30.79875, 38.36204, 47.65634, 57.61045, 69.25548, 56.99433, 
    75.02316, 89.26183, 99.31198, 105.3863, 107.4346, 105.4044, 99.39714, 
    89.63618, 76.6698, 63.14838, 86.80895, 87.42487, 90.17094,
  39.39671, 44.05953, 52.45988, 62.53069, 72.60616, 83.57346, 69.27618, 
    93.76754, 114.53, 129.5341, 138.6108, 141.6595, 138.6222, 129.596, 
    114.8998, 95.92701, 78.17574, 109.1279, 114.5359, 120.4684,
  49.38883, 53.38571, 60.33288, 67.7957, 73.53912, 77.97214, 63.23856, 
    88.99162, 113.5822, 132.4919, 144.2536, 148.2357, 144.2435, 132.4898, 
    113.9222, 91.84297, 74.99574, 109.9615, 123.7914, 134.4966,
  53.72971, 56.49231, 60.4273, 62.66714, 60.84435, 55.45491, 35.85291, 
    55.8143, 77.86352, 96.38158, 108.6471, 112.9233, 108.5966, 96.2973, 
    78.29782, 59.89732, 51.26128, 90.55229, 113.6843, 129.7415,
  48.09336, 49.69988, 50.85714, 48.78748, 41.80927, 30.98616, 10.34214, 
    21.5361, 34.74971, 46.08889, 53.906, 56.71057, 53.91137, 46.24279, 
    35.87788, 26.74474, 26.02831, 62.24679, 87.66895, 104.9323,
  33.65225, 34.37014, 33.97928, 30.62699, 23.76521, 14.57213, 0.5375938, 
    4.574684, 9.069759, 12.48733, 14.81139, 15.67383, 14.91765, 12.95355, 
    10.73814, 9.524582, 12.23051, 36.18205, 54.70992, 67.10248,
  15.95618, 15.81433, 14.71844, 12.20469, 8.613858, 4.630041, -0.424257, 
    -1.303278, -2.186762, -3.087647, -3.690042, -3.879523, -3.593663, 
    -2.719116, -1.049409, 1.616113, 5.671009, 14.92025, 22.34952, 27.04918,
  -10.57996, -11.96049, -14.03462, -15.87991, -16.8737, -17.02542, -17.02045, 
    -18.22272, -19.48336, -20.70046, -21.66051, -22.05468, -21.77781, 
    -21.08254, -20.4967, -20.54256, -21.60598, -24.93274, -28.69957, -31.2199,
  -27.15679, -30.48529, -35.65695, -40.63282, -43.93544, -45.625, -47.51319, 
    -54.54661, -61.23045, -66.88022, -70.87529, -72.39201, -71.14869, 
    -67.7861, -63.68253, -60.26037, -58.93343, -65.52555, -73.896, -79.78738,
  -43.65016, -47.26183, -53.05297, -58.97731, -63.4222, -66.52482, -69.51241, 
    -82.62701, -94.86787, -104.8146, -111.5984, -114.1218, -112.0361, 
    -106.2622, -98.77639, -91.6667, -87.27901, -96.7786, -107.6445, -115.4572,
  -58.97543, -61.36917, -65.65294, -70.65129, -74.97813, -78.73692, 
    -80.39551, -98.73148, -115.863, -129.5299, -138.6638, -142.0157, 
    -139.215, -131.384, -120.9545, -110.6275, -103.657, -117.4137, -129.4714, 
    -138.2705,
  -72.14185, -72.6461, -74.49891, -77.6414, -80.89789, -84.26846, -81.29797, 
    -103.4032, -124.6502, -141.7997, -153.2498, -157.394, -153.7365, 
    -143.5929, -130.0563, -117.0471, -109.0564, -129.8989, -143.003, -152.6527,
  -82.76282, -81.4641, -80.91291, -81.93651, -83.51402, -85.66055, -75.37763, 
    -100.0129, -125.1618, -146.3909, -160.8042, -165.9149, -160.8438, 
    -147.0778, -128.9846, -113.3884, -106.6979, -137.6616, -152.1999, 
    -162.9026,
  -86.05029, -84.03404, -82.81857, -83.74482, -85.80144, -88.87813, 
    -72.29118, -97.9371, -124.0907, -146.0482, -160.6812, -165.7679, 
    -160.5644, -146.1696, -126.555, -109.3319, -101.9986, -142.553, 
    -155.9235, -165.8168,
  -80.14867, -78.54375, -78.33862, -80.96058, -85.35819, -91.26983, 
    -72.39513, -97.04541, -120.5032, -139.0717, -150.8552, -154.8716, 
    -150.8622, -139.3234, -122.4632, -105.8287, -96.27268, -140.0555, 
    -149.8331, -157.3463,
  -67.35779, -66.47896, -67.34962, -71.14803, -76.95428, -84.62107, 
    -66.21383, -87.79704, -106.7686, -120.844, -129.4121, -132.2907, 
    -129.4591, -121.1045, -108.2263, -94.28362, -84.86259, -124.4407, 
    -130.6207, -135.7969,
  -48.58047, -48.31433, -49.67328, -53.4353, -58.93221, -66.17633, -51.53963, 
    -67.47118, -80.47068, -89.63609, -95.08163, -96.90305, -95.14078, 
    -89.88199, -81.53403, -71.83743, -64.40726, -94.12023, -97.33977, 
    -100.4465,
  -25.45975, -25.47845, -26.49236, -28.87106, -32.2582, -36.69002, -28.46123, 
    -36.83319, -43.34578, -47.81297, -50.44235, -51.32278, -50.48307, 
    -47.97033, -43.94495, -39.09209, -35.07424, -51.09943, -52.3298, -53.71973,
  -0.07858224, -0.1415867, -0.2753838, -0.4864335, -0.7547989, -0.9910976, 
    -0.52315, -0.4871296, -0.4673645, -0.4632723, -0.4683489, -0.4721751, 
    -0.4712813, -0.4751819, -0.5051452, -0.5742351, -0.6532062, -1.181325, 
    -0.993185, -0.8325638,
  25.16629, 24.97234, 25.54023, 27.22103, 29.7024, 33.23046, 26.43545, 
    34.84439, 41.42812, 45.9366, 48.57104, 49.44621, 48.59969, 46.0464, 
    41.88456, 36.80377, 32.64899, 47.11473, 49.07212, 50.98605,
  47.75345, 46.96265, 47.23743, 49.31829, 52.57285, 57.23235, 45.39106, 
    60.91175, 73.94767, 83.24213, 88.75664, 90.58734, 88.77728, 83.34618, 
    74.63119, 64.59949, 57.47618, 84.20755, 89.4758, 93.80547,
  65.21203, 63.13875, 61.57753, 61.6527, 62.43466, 63.81596, 49.30069, 
    68.20686, 86.09529, 99.90751, 108.4564, 111.3223, 108.4048, 99.84698, 
    86.83084, 73.61968, 66.76589, 101.7821, 112.7376, 120.446,
  75.259, 71.31387, 66.45077, 62.14444, 57.38316, 51.74424, 34.71607, 
    51.22237, 69.18611, 84.50061, 94.66908, 98.17429, 94.52256, 84.33943, 
    70.40363, 59.03139, 57.18952, 96.72884, 114.6009, 126.1553,
  76.26847, 70.36334, 61.67908, 52.0811, 41.0761, 28.71839, 5.972911, 
    17.75934, 31.70894, 44.13129, 52.801, 55.84736, 52.57582, 44.01205, 
    33.71798, 28.07047, 32.90111, 74.69729, 97.01473, 111.2593,
  65.44547, 58.75645, 48.36352, 36.57188, 23.72631, 10.39655, -11.20829, 
    -3.660346, 4.72131, 11.54167, 16.17674, 17.83229, 16.24694, 12.24578, 
    8.137508, 7.497114, 13.70389, 48.63504, 68.41103, 81.12988,
  45.14243, 39.50257, 30.74117, 21.21976, 11.7321, 2.644737, -10.95535, 
    -7.769814, -5.018127, -3.601294, -2.89098, -2.575095, -2.426585, 
    -2.042631, -0.7839279, 1.861667, 6.593771, 27.68835, 39.55094, 46.94751,
  21.50693, 18.24981, 13.32874, 8.425217, 4.242831, 0.7613497, -3.701637, 
    -4.468724, -5.797777, -7.521692, -8.897655, -9.322088, -8.457384, 
    -6.233342, -2.801038, 1.356099, 5.501413, 12.43878, 15.86745, 17.58074,
  -15.66589, -15.82209, -15.83138, -15.34673, -14.20648, -12.55131, 
    -10.72263, -10.16477, -9.517902, -8.877159, -8.454716, -8.383898, 
    -8.783413, -9.800936, -11.60561, -14.25838, -17.68761, -22.95474, 
    -27.73217, -30.66876,
  -38.78097, -39.26811, -39.70596, -39.33284, -37.58064, -34.73182, -31.6505, 
    -34.27618, -36.51506, -38.12688, -39.27155, -39.85835, -39.98368, 
    -40.18206, -41.30058, -43.91034, -48.37148, -60.26365, -71.44547, 
    -78.61004,
  -59.42254, -59.28409, -59.07399, -58.49114, -56.89332, -54.49013, 
    -51.00517, -58.60975, -65.50463, -70.83438, -74.50591, -76.07648, 
    -75.56312, -73.91054, -72.7151, -73.14291, -76.05782, -92.30894, 
    -106.2736, -115.3946,
  -76.44374, -74.96587, -73.23466, -71.96081, -70.6693, -69.43098, -64.80992, 
    -78.05393, -90.45532, -100.2985, -107.0143, -109.7045, -108.2537, 
    -103.9957, -99.33739, -96.27352, -96.34055, -116.4141, -130.6173, 
    -140.1768,
  -89.74647, -86.70622, -83.05086, -80.53857, -78.95724, -78.33524, 
    -70.25279, -88.15631, -105.569, -119.8134, -129.5478, -133.2559, 
    -130.5969, -123.2644, -114.7094, -108.4108, -106.7362, -132.3715, 
    -146.2096, -155.8683,
  -99.97684, -95.41449, -89.65981, -85.3273, -82.56188, -81.51907, -67.82377, 
    -88.76983, -110.304, -128.754, -141.5144, -146.0854, -141.6755, 
    -130.3433, -117.3172, -109.0121, -108.452, -141.9214, -155.7796, -165.6759,
  -102.8937, -97.73713, -91.33127, -86.76258, -84.30923, -84.02121, -65.566, 
    -87.55258, -110.2377, -129.7502, -143.0573, -147.6875, -142.8529, 
    -130.2649, -115.2127, -105.3666, -104.3441, -145.8865, -158.2497, 
    -167.1171,
  -96.4743, -91.73599, -86.24565, -83.1283, -82.57418, -84.34652, -64.39747, 
    -85.39906, -106.0414, -123.0425, -134.1307, -137.9338, -134.1122, 
    -123.5783, -109.8651, -99.40062, -96.0727, -140.7012, -150.1302, -156.9265,
  -82.1479, -78.23842, -74.01793, -72.2993, -73.23328, -76.48003, -57.5843, 
    -76.09214, -93.1859, -106.3832, -114.5524, -117.2988, -114.592, -106.798, 
    -95.84843, -86.50914, -82.5813, -122.7384, -129.2196, -133.9787,
  -60.11056, -57.34661, -54.56653, -53.91239, -55.49525, -59.00305, 
    -44.22226, -58.13086, -70.11179, -78.78861, -83.94595, -85.6621, 
    -84.01486, -79.12848, -71.85828, -65.0263, -61.5969, -91.67543, 
    -95.47868, -98.36955,
  -31.90625, -30.52489, -29.25553, -29.25474, -30.5624, -32.94227, -24.50672, 
    -31.90546, -37.96257, -42.17449, -44.62767, -45.44399, -44.68398, 
    -42.39764, -38.90644, -35.43764, -33.52331, -49.95691, -51.56145, 
    -52.81517,
  -0.3468877, -0.5316474, -0.8979084, -1.429372, -2.065024, -2.633322, 
    -1.438333, -1.351082, -1.269208, -1.21503, -1.193636, -1.192821, 
    -1.212038, -1.27977, -1.439045, -1.664361, -1.82546, -3.165782, -2.76039, 
    -2.439,
  30.81137, 28.89671, 26.57265, 25.03687, 24.45812, 24.94188, 19.66735, 
    27.07566, 33.33033, 37.74308, 40.30568, 41.13987, 40.29553, 37.74342, 
    33.73499, 29.71516, 27.67584, 40.62255, 43.58016, 45.75403,
  57.59688, 53.771, 48.89949, 45.19191, 42.8869, 41.91228, 32.0792, 44.85047, 
    56.69673, 65.66752, 71.09354, 72.86996, 70.98973, 65.48413, 57.35673, 
    50.23409, 47.89017, 72.36665, 79.29023, 83.94828,
  76.5958, 70.67654, 62.52936, 55.1106, 48.69528, 42.90662, 29.83645, 
    43.46108, 57.9833, 70.23914, 78.21806, 80.8855, 77.92639, 69.78948, 
    59.15187, 52.04794, 52.70498, 84.98363, 97.40054, 105.1716,
  85.4677, 77.44116, 65.63273, 53.55763, 41.70742, 29.7163, 13.00439, 
    23.33967, 35.92255, 47.56299, 55.74765, 58.56649, 55.37402, 47.32583, 
    38.57984, 35.68829, 41.65598, 77.82616, 95.22057, 105.8207,
  83.46524, 73.79543, 58.95757, 42.97409, 26.96475, 11.2858, -10.83011, 
    -2.462232, 7.506625, 16.41286, 22.72219, 24.87297, 22.3456, 16.53535, 
    11.47821, 12.56692, 21.59854, 58.36709, 76.93964, 88.56215,
  69.29787, 59.74027, 44.98536, 29.20876, 13.97319, -0.003744125, -20.25493, 
    -13.43172, -6.41786, -1.049319, 2.49432, 3.754521, 2.697879, 0.3533792, 
    -0.9390578, 1.43495, 8.078769, 37.44561, 51.74565, 61.00172,
  46.62874, 39.3455, 28.29105, 16.95876, 6.710728, -2.119018, -14.72488, 
    -11.35695, -8.632333, -7.27468, -6.593684, -6.180603, -5.691177, 
    -4.618644, -2.426584, 0.7805189, 4.374966, 21.30733, 28.7139, 33.42551,
  21.96922, 18.22224, 12.65127, 7.261942, 2.876321, -0.5538176, -4.759269, 
    -5.359424, -6.488529, -7.983994, -9.13667, -9.353234, -8.257927, 
    -5.718797, -1.975113, 2.079956, 5.162745, 9.969095, 11.34489, 11.92048,
  -21.5704, -19.71292, -16.63556, -13.11727, -9.62239, -6.310662, -2.955809, 
    -1.084725, 0.9087341, 2.782294, 4.025656, 4.209105, 3.047553, 0.4450922, 
    -3.429473, -8.011736, -12.51023, -17.86747, -21.63941, -23.70904,
  -51.77546, -47.79446, -41.2298, -33.6713, -25.94962, -18.51899, -10.69892, 
    -9.526765, -8.043713, -6.370691, -5.336001, -5.495491, -7.31543, 
    -11.24329, -17.42186, -25.06025, -32.88824, -46.63835, -56.70504, 
    -62.70368,
  -76.88577, -71.51176, -62.83322, -53.06315, -43.19859, -33.82847, 
    -22.64277, -23.98984, -24.90462, -25.14243, -25.50576, -26.38068, 
    -28.27309, -32.05412, -38.41264, -46.67517, -55.43565, -75.89024, 
    -89.74456, -98.26817,
  -95.82471, -89.67996, -80.01942, -69.52985, -59.31784, -50.08677, 
    -36.34429, -42.02641, -47.35846, -51.41029, -54.47461, -56.39481, 
    -57.54406, -59.31385, -63.31595, -69.61649, -77.07286, -102.7289, 
    -117.6539, -127.1955,
  -109.2297, -102.5367, -92.23365, -81.41008, -71.39154, -63.11453, 
    -46.68382, -57.12807, -67.63763, -76.39143, -82.73289, -85.66451, 
    -85.2968, -83.6619, -83.79886, -87.26824, -93.17207, -123.5026, -137.764, 
    -147.3091,
  -118.3712, -110.9597, -99.59579, -87.81447, -77.40036, -69.64233, 
    -50.31886, -64.34573, -79.28471, -92.35977, -101.6509, -105.1009, 
    -102.4635, -96.67115, -93.0112, -95.19656, -101.6147, -136.2736, 
    -149.2892, -158.3145,
  -119.6275, -112.0846, -100.6217, -88.95564, -79.0207, -72.06384, -51.27093, 
    -66.91423, -83.72282, -98.69751, -109.2257, -112.838, -109.0594, 
    -100.852, -94.44549, -94.88575, -100.4824, -139.5073, -150.526, -158.1837,
  -111.1488, -104.2501, -93.97078, -83.87133, -75.66946, -70.2076, -49.73266, 
    -64.88419, -80.83105, -94.90045, -104.5628, -107.8829, -104.4914, 
    -96.44669, -89.01405, -87.29229, -90.4179, -131.3437, -139.8648, -145.6557,
  -94.06003, -88.2375, -79.69209, -71.56972, -65.33984, -61.49834, -42.77941, 
    -56.19501, -70.00492, -81.69579, -89.32969, -91.88576, -89.24643, 
    -82.56604, -75.66946, -73.26839, -75.14549, -111.7154, -117.7993, 
    -121.8099,
  -68.66805, -64.47958, -58.42404, -52.87185, -48.90326, -46.71387, 
    -32.08043, -42.37986, -52.57434, -60.6961, -65.71739, -67.36491, 
    -65.68513, -61.17919, -56.06732, -53.86819, -54.88831, -82.46386, 
    -86.22298, -88.60812,
  -36.83711, -34.82021, -32.0102, -29.64484, -28.23645, -27.71481, -18.59245, 
    -24.139, -29.4097, -33.39837, -35.77774, -36.56231, -35.8253, -33.76416, 
    -31.33343, -30.26199, -30.80379, -46.85652, -48.39365, -49.29544,
  -1.878941, -2.454719, -3.540194, -5.012104, -6.690383, -8.27239, -4.79596, 
    -4.646171, -4.343847, -4.037084, -3.849496, -3.826527, -4.017534, 
    -4.510039, -5.25757, -5.878612, -6.044298, -10.04886, -9.172229, -8.555359,
  31.82194, 28.40066, 22.93327, 16.92274, 11.22472, 6.256028, 4.940283, 
    10.04394, 15.67746, 20.36023, 23.25811, 24.10953, 22.80649, 19.42477, 
    15.33218, 13.37345, 14.36884, 21.18471, 25.17556, 27.59805,
  59.62546, 53.33162, 43.27343, 32.13936, 21.30409, 11.11545, 5.769981, 
    12.6843, 21.49644, 29.64604, 35.09272, 36.72816, 34.17775, 28.13339, 
    22.053, 20.92716, 25.03065, 40.30295, 48.33565, 52.95118,
  77.65317, 68.80677, 54.50928, 38.31799, 21.99139, 5.888213, -3.632551, 
    1.283457, 9.253246, 17.66452, 23.84552, 25.75103, 22.75389, 16.5553, 
    12.25319, 15.01645, 23.65347, 44.52274, 56.58503, 63.40143,
  83.7362, 73.16293, 55.90674, 36.07452, 15.8522, -3.880921, -17.93824, 
    -14.86372, -9.171947, -2.951855, 1.855091, 3.375387, 1.178333, -2.581316, 
    -3.128782, 3.180562, 14.21863, 37.5198, 51.36851, 59.45562,
  78.26124, 67.26434, 49.20829, 28.42206, 7.592715, -11.50933, -30.37125, 
    -25.09928, -18.72429, -13.22434, -9.403397, -8.267683, -9.832298, 
    -12.12834, -11.49871, -5.560964, 3.404448, 26.72626, 38.65306, 46.33313,
  61.93703, 52.63033, 37.36197, 19.94074, 2.921275, -11.79799, -29.17885, 
    -23.02537, -16.91024, -12.42624, -9.551826, -8.499173, -9.004934, 
    -9.780152, -8.929657, -5.699396, -1.870447, 16.82608, 24.39277, 29.91615,
  39.8352, 33.86643, 24.04607, 12.89303, 2.162411, -6.893585, -18.13376, 
    -14.65759, -11.59925, -9.6921, -8.46126, -7.601556, -6.751884, -5.421879, 
    -3.444169, -1.624075, -1.195915, 9.451502, 12.68241, 15.32838,
  18.20193, 15.83137, 11.72931, 6.898303, 2.241995, -1.671676, -5.855297, 
    -6.347271, -6.932801, -7.623755, -7.988453, -7.619825, -6.214831, 
    -3.726157, -0.674961, 1.749157, 2.512173, 4.744701, 4.806832, 4.964711,
  -22.78646, -20.32372, -16.26666, -11.694, -7.29075, -3.316508, 0.5938988, 
    2.742913, 4.832452, 6.644944, 7.705643, 7.614685, 6.107108, 3.136334, 
    -0.9762162, -5.410746, -9.188211, -13.49923, -16.05621, -17.39629,
  -54.37465, -48.88456, -39.82329, -29.504, -19.35097, -10.10894, -0.5062761, 
    1.697052, 3.894907, 5.963169, 7.038784, 6.513466, 3.902041, -1.11741, 
    -8.280678, -16.16011, -22.98361, -35.20954, -42.90702, -47.46625,
  -80.91904, -73.67202, -61.66471, -47.8269, -33.95269, -21.18949, -6.493052, 
    -5.361341, -4.234306, -2.996913, -2.639496, -3.753462, -6.935965, 
    -12.84844, -21.51448, -31.30702, -40.04369, -59.83308, -71.56388, 
    -78.78355,
  -101.11, -93.20427, -80.1215, -64.95736, -49.60473, -35.54214, -16.75195, 
    -18.28936, -19.96803, -21.18319, -22.60651, -24.4651, -27.32714, -32.34, 
    -40.25465, -49.91657, -59.0913, -85.4659, -99.30655, -108.138,
  -115.0628, -106.9831, -93.69126, -78.32533, -62.86846, -49.12922, 
    -27.35186, -32.58488, -38.38119, -43.37324, -47.39198, -49.93434, 
    -51.43685, -53.7994, -59.12725, -67.43405, -76.34633, -107.714, 
    -121.6206, -130.8412,
  -123.6131, -115.2809, -101.616, -85.90762, -70.46558, -57.46745, -34.22916, 
    -42.70699, -52.60939, -61.549, -68.09686, -70.7815, -69.94392, -68.72716, 
    -71.33198, -79.12908, -88.69624, -122.6311, -135.2538, -143.8687,
  -123.4817, -115.4434, -102.3341, -87.36015, -72.80404, -60.76189, 
    -38.46811, -49.04274, -61.44747, -72.92484, -81.15329, -83.96485, 
    -81.43056, -77.18964, -76.79473, -82.68567, -91.2338, -126.707, 
    -137.3206, -144.5293,
  -113.3639, -106.2933, -94.88679, -81.9927, -69.48563, -58.98208, -38.48302, 
    -49.37969, -61.97391, -73.7709, -82.1842, -85.04858, -82.19771, -76.6199, 
    -73.74438, -76.60625, -82.46851, -118.703, -126.9852, -132.4395,
  -94.86278, -89.11125, -79.90287, -69.59222, -59.66298, -51.2742, -32.77839, 
    -42.55191, -53.91412, -64.36797, -71.53465, -73.89072, -71.33763, 
    -65.94521, -62.31736, -63.6816, -67.91669, -100.4127, -106.3555, -110.1124,
  -68.91152, -64.95608, -58.68034, -51.74071, -45.13377, -39.51592, -24.6404, 
    -32.20193, -40.91321, -48.56927, -53.54359, -55.1332, -53.36432, 
    -49.3693, -46.28081, -46.84621, -49.7169, -74.84649, -78.54544, -80.74909,
  -37.69104, -36.00185, -33.42338, -30.72431, -28.29621, -26.26653, 
    -15.92116, -19.98517, -24.51894, -28.29597, -30.64993, -31.42566, 
    -30.71591, -29.01246, -27.73923, -28.23662, -29.79964, -45.90371, 
    -47.329, -48.07955,
  -4.484623, -5.44755, -7.23865, -9.62833, -12.34484, -15.04646, -9.118135, 
    -9.098068, -8.625631, -8.008554, -7.589539, -7.578354, -8.129895, 
    -9.296906, -10.64974, -11.39457, -11.31205, -18.50602, -17.31887, 
    -16.55667,
  26.60155, 22.75922, 16.15751, 8.021649, -0.7744622, -9.626503, -7.660074, 
    -4.949342, -0.2908468, 4.455471, 7.653962, 8.397605, 6.35127, 2.168941, 
    -1.385203, -1.374341, 1.516347, 1.893377, 6.323151, 8.805396,
  51.35007, 44.6983, 33.34238, 19.38106, 4.153732, -11.644, -13.76837, 
    -11.65632, -6.004647, 0.6540661, 5.562976, 6.745186, 3.642213, -1.874174, 
    -4.886171, -1.725531, 5.397996, 11.52582, 19.5729, 23.91273,
  66.43714, 57.54219, 42.35634, 23.6286, 3.098215, -18.22609, -24.95571, 
    -25.2482, -21.65744, -16.39505, -12.0913, -11.02792, -13.63849, 
    -17.24487, -16.71908, -9.45707, 1.250368, 11.22685, 22.01423, 27.90869,
  70.41347, 60.43116, 43.36805, 22.31733, -0.5501938, -23.4579, -34.87513, 
    -35.06982, -32.48489, -28.93202, -25.9916, -25.19734, -26.55371, 
    -27.5827, -24.49831, -16.04114, -5.492265, 6.511325, 17.54491, 24.03288,
  64.40004, 54.77932, 38.26867, 17.94546, -3.610199, -23.75947, -39.78115, 
    -36.11964, -31.18216, -26.98171, -24.17397, -23.44648, -24.44451, 
    -25.11479, -22.76836, -16.78775, -10.09875, 3.079167, 11.40567, 17.16373,
  49.68702, 42.27765, 29.44221, 13.54367, -3.13631, -17.98916, -33.34951, 
    -28.1025, -22.57471, -18.46113, -15.83461, -14.83864, -15.07872, 
    -15.32297, -14.28725, -12.06656, -10.5884, 1.188962, 5.864606, 9.917366,
  31.08326, 26.95424, 19.54571, 9.994987, -0.3009566, -9.523952, -19.95809, 
    -16.85095, -13.81059, -11.6366, -10.06671, -8.932133, -7.975448, 
    -6.902313, -5.838289, -5.597525, -7.014921, 0.1256447, 1.98228, 4.051605,
  13.8562, 12.73114, 10.26664, 6.495584, 2.026681, -2.193106, -6.431762, 
    -6.993981, -7.288335, -7.451492, -7.259804, -6.473562, -4.946119, 
    -2.852499, -0.9026124, -0.04551804, -0.6194304, 0.5310047, 0.4533701, 
    0.7020123,
  -21.47739, -19.18572, -15.24336, -10.52808, -5.74851, -1.367111, 2.889592, 
    5.063458, 6.908729, 8.293149, 8.875579, 8.381845, 6.656716, 3.773781, 
    0.1889415, -3.228668, -5.666788, -8.762212, -10.33499, -11.19886,
  -51.4446, -45.97021, -36.66043, -25.60985, -14.38914, -4.157184, 6.48876, 
    9.03833, 11.14736, 12.79068, 13.26795, 12.11983, 9.02669, 3.924657, 
    -2.570264, -8.808918, -13.17458, -23.12204, -28.51875, -31.88545,
  -77.77494, -70.22198, -57.32809, -41.82443, -25.75718, -10.8723, 6.039184, 
    8.524315, 10.43647, 11.90846, 12.03847, 10.31194, 6.294738, -0.2942963, 
    -8.912996, -17.53048, -23.97034, -41.44839, -50.50821, -56.30569,
  -98.78069, -90.26899, -75.69456, -57.93658, -39.16296, -21.54646, 
    0.8166075, 2.281775, 2.978539, 3.346961, 2.605844, 0.4091721, -3.742411, 
    -10.53003, -19.89841, -30.00835, -38.31121, -63.16307, -74.92683, 
    -82.61201,
  -113.5045, -104.7602, -89.79615, -71.43068, -51.83174, -33.4715, -7.443206, 
    -7.988832, -9.736576, -11.65077, -13.89711, -16.35942, -19.60811, 
    -25.06937, -33.73888, -44.48233, -54.26244, -84.60802, -97.37608, 
    -105.8955,
  -121.8835, -113.1379, -98.18414, -79.80933, -60.33012, -42.46923, 
    -15.80936, -18.44718, -23.23953, -28.1018, -32.02351, -34.20916, 
    -35.51253, -38.70344, -46.33142, -57.87823, -69.22669, -101.1025, 
    -113.1905, -121.3536,
  -120.8873, -112.8214, -99.04983, -82.0502, -63.87702, -47.02449, -23.36041, 
    -28.19664, -35.76738, -43.42666, -49.10954, -51.21132, -50.50024, 
    -50.67891, -55.67075, -65.6675, -76.37912, -107.288, -117.8423, -124.8266,
  -109.8819, -103.1312, -91.65424, -77.39805, -61.7991, -46.73886, -26.31367, 
    -32.51496, -41.43057, -50.6004, -57.41776, -59.73906, -57.86215, 
    -55.38795, -56.86255, -63.30333, -71.24992, -101.8032, -110.2997, 
    -115.7166,
  -91.16029, -85.96675, -77.16202, -66.16157, -53.90265, -41.70652, 
    -23.29541, -29.17344, -37.78896, -46.66543, -53.0885, -55.13578, 
    -52.94581, -49.514, -49.24625, -53.54484, -59.44482, -87.42096, 
    -93.55708, -97.32095,
  -66.38305, -63.06902, -57.48158, -50.46671, -42.49192, -34.26954, 
    -18.62589, -23.20691, -30.07144, -36.95935, -41.72374, -43.18835, 
    -41.49056, -38.60871, -37.91448, -40.73537, -44.84127, -67.78362, 
    -71.60989, -73.8224,
  -38.01566, -36.90614, -35.12104, -32.91761, -30.33075, -27.48783, 
    -15.15728, -17.63836, -21.1812, -24.53911, -26.77251, -27.54697, 
    -27.05267, -26.17779, -26.39146, -28.1563, -30.28642, -47.35542, 
    -48.76654, -49.49801,
  -9.160686, -10.52191, -13.04525, -16.41547, -20.31723, -24.46612, 
    -15.52223, -16.02203, -15.57669, -14.67111, -14.00553, -14.13589, 
    -15.35538, -17.38744, -19.11898, -19.58108, -18.98727, -30.73553, 
    -29.34264, -28.54416,
  16.65107, 12.71881, 5.676953, -3.63409, -14.65905, -26.94499, -21.65279, 
    -22.12616, -19.33148, -15.2029, -12.12229, -11.81321, -14.68689, 
    -18.93054, -20.81589, -18.50838, -13.99399, -21.55243, -16.93452, 
    -14.51383,
  36.11775, 29.85812, 18.71854, 3.982921, -13.60238, -33.4165, -32.46523, 
    -35.24529, -33.39664, -29.17287, -25.6356, -25.26806, -28.36839, 
    -31.87978, -31.08309, -24.6434, -15.94534, -20.27914, -12.63268, -8.665838,
  47.1015, 39.25946, 25.33849, 6.928623, -14.95528, -39.13197, -42.89997, 
    -47.31739, -47.41232, -45.10374, -42.80022, -42.54561, -44.25959, 
    -44.95516, -40.94123, -31.87442, -21.34969, -23.07173, -13.76743, 
    -8.702431,
  49.32507, 41.08102, 26.44262, 7.100397, -15.56757, -39.48875, -47.87655, 
    -50.40115, -49.932, -48.20572, -46.60143, -46.24586, -46.75249, 
    -45.90194, -41.39438, -33.40509, -24.90522, -24.19529, -15.51314, 
    -10.20737,
  44.47781, 37.01419, 23.69954, 6.124193, -13.96864, -33.75528, -46.63371, 
    -44.72972, -41.05537, -37.81411, -35.73158, -35.25153, -35.77156, 
    -35.52611, -32.93655, -28.2904, -24.04869, -20.32892, -14.56847, -10.12261,
  33.63022, 28.30291, 18.63852, 5.625404, -9.290783, -23.45269, -36.58985, 
    -32.79657, -28.18752, -24.59452, -22.29, -21.3996, -21.49671, -21.60775, 
    -21.04398, -20.17264, -20.44373, -14.83411, -12.04777, -8.977339,
  20.44341, 17.88276, 12.91302, 5.605396, -3.377453, -12.21528, -21.65387, 
    -19.26658, -16.59128, -14.43278, -12.73302, -11.49199, -10.63996, 
    -10.13679, -10.23746, -11.41141, -13.95165, -9.803828, -8.758239, 
    -7.067507,
  8.923646, 8.652339, 7.586374, 5.142548, 1.40625, -2.695833, -6.810647, 
    -7.527549, -7.693503, -7.487506, -6.859431, -5.770658, -4.321906, 
    -2.942648, -2.322141, -2.863278, -4.276811, -3.873793, -3.958372, 
    -3.641281,
  -16.0425, -14.7306, -12.17116, -8.540133, -4.232083, 0.1008631, 4.448836, 
    6.429172, 7.744714, 8.362329, 8.169736, 7.162766, 5.47149, 3.418932, 
    1.514658, 0.2985373, -0.02675784, -1.640656, -2.312912, -2.8362,
  -39.00587, -35.20025, -28.28275, -19.15114, -8.811997, 1.260757, 12.27288, 
    14.72568, 16.22031, 16.81637, 16.16279, 14.23262, 11.20504, 7.504007, 
    3.936111, 1.690735, 1.46381, -5.30113, -8.186871, -10.41326,
  -61.17845, -55.18677, -44.49855, -30.61987, -14.98501, 0.3070831, 18.19406, 
    21.31667, 23.18855, 23.93972, 23.03439, 20.44182, 16.34989, 11.15456, 
    5.74538, 1.723902, 0.3582659, -12.66139, -18.02501, -22.01751,
  -80.92233, -73.32594, -59.8993, -42.55385, -22.94476, -3.556789, 20.7704, 
    24.59884, 26.83661, 27.73166, 26.71965, 23.80584, 19.10056, 12.76098, 
    5.456597, -1.109735, -4.983278, -24.8284, -32.65542, -38.29974,
  -96.09644, -87.66845, -72.82404, -53.62873, -31.80178, -9.990019, 18.87824, 
    23.31131, 25.57882, 26.27139, 25.13446, 22.27239, 17.54366, 10.56056, 
    1.46416, -8.155136, -15.5037, -40.77286, -50.4795, -57.29284,
  -105.2381, -96.6762, -81.58575, -61.99783, -39.65856, -17.20201, 12.09322, 
    17.27609, 19.15248, 19.1394, 17.87403, 15.5485, 11.34643, 3.93097, 
    -7.117217, -20.08755, -31.21833, -57.31314, -67.79276, -74.90237,
  -105.2552, -97.57866, -83.98596, -66.05049, -45.0244, -23.01504, 1.733716, 
    5.981105, 6.171741, 4.39635, 2.309849, 0.522583, -2.256998, -8.381555, 
    -19.00495, -32.5673, -45.16247, -67.82597, -78.38455, -85.11723,
  -95.97137, -89.91541, -79.14777, -64.59, -46.68755, -26.69556, -6.628879, 
    -4.890242, -7.192011, -11.4016, -15.08528, -16.75214, -17.50226, 
    -20.42348, -27.64028, -38.23794, -48.88999, -70.07344, -79.51178, 
    -85.22105,
  -80.34577, -76.09423, -68.51663, -58.02795, -44.54586, -28.68732, 
    -10.21891, -9.683882, -13.15548, -18.55935, -22.9873, -24.5011, 
    -23.98944, -24.76614, -29.36695, -37.15587, -45.19662, -66.57883, 
    -73.63666, -77.79156,
  -60.87581, -58.55809, -54.43494, -48.54198, -40.5032, -30.44833, -12.94695, 
    -12.84457, -16.01701, -20.75344, -24.51993, -25.75546, -25.14977, 
    -25.35221, -28.41831, -33.77965, -39.20061, -60.30119, -64.73881, 
    -67.27587,
  -40.31931, -40.01347, -39.52835, -38.66402, -37.01399, -34.49392, 
    -18.37363, -18.86355, -20.60171, -22.85202, -24.64096, -25.59648, 
    -26.19428, -27.40987, -29.69494, -32.4673, -34.83006, -55.64042, 
    -57.27898, -58.22304,
  -21.35233, -23.04008, -26.20275, -30.55357, -35.91483, -42.3496, -28.65363, 
    -31.11493, -31.80909, -31.27762, -30.82114, -31.66613, -33.97666, 
    -36.43351, -37.41665, -36.62444, -35.00271, -55.89157, -54.43112, 
    -53.77441,
  -6.269605, -9.732304, -16.16583, -25.31288, -37.35112, -52.59797, 
    -42.59423, -48.57256, -50.35238, -49.19701, -47.91777, -48.7968, 
    -51.56752, -53.27554, -51.33877, -46.17722, -40.24559, -61.15063, 
    -56.6156, -54.41476,
  3.628115, -1.109106, -9.894537, -22.56001, -39.5359, -61.0173, -55.37908, 
    -64.14362, -68.02122, -68.33722, -67.84585, -68.60985, -70.05829, 
    -69.33401, -64.40819, -56.21559, -47.62134, -67.68943, -60.90344, 
    -57.41985,
  8.522066, 3.234844, -6.557065, -20.77483, -39.83711, -63.28061, -61.93872, 
    -70.24364, -74.34054, -75.46165, -75.54418, -75.8782, -75.91908, 
    -73.81142, -68.38091, -60.4418, -52.34424, -70.12724, -62.64748, -58.40075,
  9.776542, 4.685036, -4.715266, -18.37911, -36.48001, -57.75269, -60.67841, 
    -65.56693, -67.36455, -67.4603, -67.08579, -66.95177, -66.64085, 
    -65.04538, -61.45629, -56.29064, -51.14726, -64.87561, -58.53009, 
    -54.30035,
  9.051078, 4.667328, -3.356376, -14.87833, -29.67484, -45.96892, -53.18661, 
    -54.31901, -52.90706, -51.11596, -49.9524, -49.70434, -49.81345, 
    -49.35739, -47.85003, -45.56541, -43.76432, -51.7372, -48.34121, -45.16394,
  6.171902, 3.218016, -2.184127, -10.05997, -20.28203, -31.31354, -40.11093, 
    -39.14405, -36.6473, -34.3303, -32.80299, -32.25876, -32.42519, 
    -32.84798, -33.31046, -33.89045, -35.24055, -37.35049, -36.31403, 
    -34.31049,
  2.802126, 1.613572, -0.6821289, -4.510668, -10.19613, -16.87631, -23.86113, 
    -22.81435, -21.22581, -19.66073, -18.27766, -17.34711, -17.11005, 
    -17.74652, -19.31893, -21.64678, -24.58378, -24.30269, -24.09835, 
    -22.96141,
  1.259096, 1.438655, 1.524176, 0.9114634, -0.9015253, -3.692018, -6.880589, 
    -7.767304, -8.010594, -7.631944, -6.746647, -5.662486, -4.874679, 
    -4.926554, -6.018282, -7.771025, -9.601748, -10.09708, -10.33669, 
    -10.13501,
  -11.21376, -10.50298, -8.970781, -6.477121, -3.109531, 0.6004732, 4.596798, 
    6.308225, 7.308775, 7.549956, 7.032943, 5.942211, 4.60816, 3.449784, 
    2.842378, 2.973505, 3.711324, 2.793286, 2.521731, 2.160635,
  -27.64134, -25.08068, -20.26864, -13.45059, -5.036229, 3.733188, 14.0797, 
    16.16479, 17.25867, 17.33427, 16.22777, 14.23675, 11.89334, 9.810631, 
    8.60747, 8.899343, 10.82026, 5.689385, 3.951624, 2.25019,
  -44.63397, -40.16193, -32.04278, -20.99927, -7.750111, 5.912923, 22.85893, 
    25.70703, 27.2515, 27.46886, 26.05779, 23.40606, 20.17022, 17.023, 
    14.66954, 14.04566, 15.74979, 5.506597, 2.066217, -0.993392,
  -61.22247, -55.01222, -43.92908, -29.17158, -11.72321, 6.279, 29.561, 
    33.67884, 36.05839, 36.7135, 35.30944, 32.29814, 28.33344, 23.95332, 
    19.73829, 16.79684, 16.42775, 0.5250807, -4.828031, -9.207532,
  -75.46683, -68.05212, -54.9071, -37.5456, -17.1211, 4.11533, 32.08504, 
    38.10869, 41.65278, 42.91422, 41.77073, 38.70392, 34.16441, 28.3274, 
    21.48087, 14.83457, 10.58117, -9.893254, -17.17738, -22.6828,
  -85.51124, -77.63484, -63.66587, -45.19907, -23.45163, -0.5397205, 
    28.11386, 36.89577, 41.93437, 43.86541, 43.23198, 40.40174, 35.23175, 
    27.36743, 16.97208, 5.594865, -3.684384, -24.4923, -33.34174, -39.48952,
  -87.98325, -80.7933, -67.94855, -50.63127, -29.55845, -6.185075, 18.09751, 
    27.66286, 32.71172, 34.33817, 33.83586, 31.5653, 26.71785, 18.25377, 
    6.12468, -7.95743, -20.69149, -37.29427, -47.55152, -53.9772,
  -82.35045, -76.72072, -66.58276, -52.48698, -34.34441, -12.66237, 6.894323, 
    14.05976, 16.84059, 16.52863, 15.08157, 13.38026, 10.31924, 4.016173, 
    -6.19578, -18.87897, -31.08947, -46.04048, -56.20556, -62.15153,
  -71.41696, -67.61391, -60.74094, -50.90126, -37.54617, -20.58609, 
    -2.096275, 2.879986, 3.727301, 1.654416, -0.8074512, -2.226466, 
    -3.794358, -7.927583, -15.59649, -25.47957, -35.01281, -52.51224, 
    -60.45952, -65.00689,
  -57.83409, -55.93701, -52.52483, -47.43444, -39.99586, -29.89625, 
    -11.16335, -8.217844, -8.351679, -10.79286, -13.32289, -14.62612, 
    -15.70468, -18.5992, -23.96702, -30.65459, -36.86199, -57.83228, 
    -62.87622, -65.7542,
  -44.33948, -44.27685, -44.2395, -43.99281, -43.09418, -41.43993, -22.99776, 
    -22.9373, -23.69343, -25.12217, -26.59551, -27.94792, -29.67595, 
    -32.19952, -35.22694, -38.12362, -40.42531, -64.98787, -66.8585, -68.02457,
  -33.14938, -34.69648, -37.65741, -41.91179, -47.53136, -54.97102, 
    -38.48101, -42.90628, -45.39814, -46.20268, -46.7029, -48.19516, 
    -50.46882, -52.00118, -51.73609, -49.99027, -47.80206, -75.48067, 
    -74.02383, -73.4893,
  -25.52044, -28.27635, -33.50854, -41.33305, -52.41468, -67.6787, -54.63039, 
    -63.68947, -69.0268, -70.92089, -71.67883, -73.0954, -74.48984, 
    -73.69647, -69.77885, -63.82951, -57.77832, -87.2048, -82.77261, -80.67523,
  -21.32314, -24.7589, -31.26222, -41.19683, -55.63335, -75.43256, -66.25295, 
    -77.27679, -84.23003, -87.36629, -88.72168, -89.68417, -89.64428, 
    -87.06636, -81.44482, -73.88265, -66.32772, -95.38107, -89.0612, -85.75684,
  -19.14935, -22.74723, -29.50538, -39.92057, -55.12923, -75.42078, 
    -69.97966, -79.3428, -85.21877, -87.97311, -89.0556, -89.42014, 
    -88.81432, -86.44443, -81.92231, -75.78252, -69.46073, -95.67999, 
    -89.01268, -85.08023,
  -17.25756, -20.62507, -26.83403, -36.31708, -49.96968, -67.43768, -65.9351, 
    -71.72894, -74.79523, -75.89434, -76.0875, -76.05216, -75.73122, 
    -74.68554, -72.48657, -69.1181, -65.46638, -86.45045, -81.06806, -77.30373,
  -14.57819, -17.49742, -22.6878, -30.29089, -40.72681, -53.25368, -55.90492, 
    -58.98654, -59.41199, -58.78931, -58.23915, -58.11998, -58.16742, 
    -57.97875, -57.27241, -55.96247, -54.76125, -68.65908, -66.22629, -63.6614,
  -12.07328, -14.03569, -17.38724, -22.21103, -28.85294, -36.74603, -41.8306, 
    -42.70027, -41.93466, -40.76233, -39.9153, -39.68495, -39.99795, 
    -40.67809, -41.55347, -42.43066, -43.66798, -49.9071, -49.61348, -48.17867,
  -8.954374, -9.692747, -10.89113, -12.82342, -16.06496, -20.50363, 
    -25.08555, -24.7627, -24.03214, -23.14175, -22.28602, -21.85655, 
    -22.20705, -23.49267, -25.55859, -27.9869, -30.61455, -32.55362, 
    -32.78402, -32.01486,
  -3.691635, -3.502691, -3.139242, -2.911201, -3.351398, -4.716835, 
    -6.696541, -7.43366, -7.758539, -7.490241, -6.776225, -6.09923, 
    -6.055148, -6.994421, -8.736481, -10.71703, -12.49206, -13.52987, 
    -13.95989, -13.9227,
  -6.092278, -5.771522, -5.037478, -3.672693, -1.535462, 1.112375, 4.364682, 
    5.638633, 6.353567, 6.388634, 5.804957, 4.931849, 4.222838, 4.06504, 
    4.605897, 5.741561, 7.1922, 6.805383, 6.884247, 6.702801,
  -15.37484, -13.76931, -10.77861, -6.359635, -0.4395463, 6.219577, 15.11567, 
    16.50376, 17.21082, 17.0324, 15.90224, 14.3636, 13.16604, 12.8987, 
    13.83226, 16.07243, 19.44951, 15.61369, 14.76845, 13.5242,
  -26.00269, -22.92129, -17.37094, -9.608732, 0.2809103, 11.09997, 25.90003, 
    27.90689, 28.99503, 28.89307, 27.43951, 25.35821, 23.61539, 22.8955, 
    23.49924, 25.71494, 29.69592, 21.8171, 19.86492, 17.57012,
  -37.88487, -33.24477, -25.00488, -13.8129, 0.0163064, 14.97205, 35.55351, 
    39.0296, 41.0938, 41.45575, 39.95676, 37.46392, 35.0426, 33.32484, 
    32.51776, 33.05382, 35.67301, 23.46166, 20.13445, 16.81462,
  -49.97295, -43.99374, -33.42466, -19.26586, -2.054826, 16.5932, 41.66457, 
    47.89623, 51.80133, 53.11935, 51.88712, 49.07139, 45.68373, 42.15935, 
    38.53928, 35.42766, 34.37299, 18.8378, 13.78026, 9.477135,
  -60.70842, -53.94305, -41.96528, -25.96003, -6.588194, 14.73369, 40.85111, 
    51.51456, 58.48825, 61.42827, 60.83582, 57.64373, 52.59534, 45.95424, 
    37.83781, 29.25177, 22.52445, 7.398888, 0.3350887, -4.790882,
  -66.57765, -60.11045, -48.55005, -32.78637, -13.06688, 9.895004, 32.59689, 
    46.00597, 54.95802, 59.10273, 59.31455, 56.30177, 50.27828, 41.21658, 
    29.38305, 16.16301, 4.212794, -6.3959, -16.01435, -21.98218,
  -66.31979, -61.12185, -51.73301, -38.50409, -20.97334, 1.093421, 19.88739, 
    31.81179, 39.59064, 43.09734, 43.45784, 41.26761, 36.10059, 27.3532, 
    15.22724, 1.249817, -12.04642, -21.28489, -31.99496, -38.08493,
  -62.02942, -58.50836, -52.13469, -42.90775, -30.03164, -12.79154, 5.65886, 
    14.76894, 20.37907, 22.297, 21.99039, 20.20809, 16.10457, 8.712366, 
    -1.669745, -13.44665, -24.46478, -38.64868, -47.50549, -52.43641,
  -55.999, -54.2509, -51.13231, -46.49342, -39.61349, -29.91, -10.28239, 
    -5.081291, -2.064192, -1.654675, -2.65672, -4.402774, -7.688489, 
    -13.24776, -20.58685, -28.43701, -35.44205, -56.83648, -62.4952, -65.71262,
  -50.57492, -50.42592, -50.28175, -50.05048, -49.45945, -48.57372, -28.4268, 
    -28.5498, -28.91562, -29.83746, -31.2009, -33.09012, -35.75926, 
    -39.01199, -42.27563, -45.13809, -47.37553, -75.90415, -77.92915, 
    -79.27623,
  -47.25802, -48.33884, -50.50392, -53.89317, -58.92099, -66.50152, 
    -47.68785, -54.01271, -58.80884, -61.74316, -63.69784, -65.53989, 
    -66.96112, -67.08775, -65.70002, -63.39091, -60.92011, -94.86034, 
    -93.31274, -92.82359,
  -46.20873, -48.05255, -51.64623, -57.43758, -66.51933, -80.3606, -64.24531, 
    -75.1257, -83.49831, -88.45677, -91.13953, -92.5619, -92.35094, 
    -89.81024, -85.13283, -79.35344, -73.68272, -110.2652, -105.8494, 
    -103.7649,
  -46.19802, -48.38004, -52.5569, -59.41321, -70.45887, -87.13258, -74.03162, 
    -85.72243, -94.71706, -100.0416, -102.6753, -103.5329, -102.5881, 
    -99.55233, -94.54167, -88.27481, -81.91293, -117.9825, -111.9809, 
    -108.7665,
  -45.29652, -47.53732, -51.69228, -58.47859, -69.43948, -85.54836, 
    -75.53341, -84.84727, -91.80791, -95.76675, -97.52103, -97.95282, 
    -97.37778, -95.67968, -92.56593, -88.09086, -83.09698, -115.6014, 
    -109.5117, -105.813,
  -42.02843, -44.16418, -47.91963, -53.80264, -63.05221, -76.12508, 
    -69.71951, -75.835, -79.95338, -82.00792, -82.74822, -82.95847, 
    -83.01541, -82.81545, -81.82019, -79.60954, -76.70949, -103.0402, 
    -98.34802, -94.971,
  -36.03347, -37.95248, -41.06981, -45.47671, -51.85477, -60.3245, -58.02722, 
    -62.64536, -64.97668, -65.64626, -65.69827, -65.68025, -65.73323, 
    -65.79404, -65.53505, -64.57446, -63.34645, -81.74197, -79.9695, -77.90598,
  -28.73282, -30.02653, -31.91583, -34.33338, -37.75725, -42.35653, 
    -43.35835, -45.67962, -46.64293, -46.70416, -46.55175, -46.59633, 
    -47.0022, -47.78056, -48.71143, -49.42986, -50.15817, -59.71394, 
    -59.91144, -58.93586,
  -19.79081, -20.24242, -20.70684, -21.22163, -22.33382, -24.423, -26.22143, 
    -26.302, -26.31841, -26.17573, -25.99826, -26.18512, -27.08599, 
    -28.76178, -30.91719, -33.08383, -35.17171, -38.99792, -39.53963, 
    -39.08194,
  -8.232371, -8.067978, -7.588739, -6.834081, -6.173195, -6.078461, 
    -6.534873, -6.805529, -7.089983, -7.048265, -6.783099, -6.790634, 
    -7.546387, -9.112827, -11.1076, -13.0327, -14.64354, -16.15978, 
    -16.76531, -16.88326,
  1.395123, 1.411376, 1.387794, 1.40718, 1.696909, 2.360362, 3.908303, 
    4.130847, 4.346314, 4.340132, 4.152769, 4.131593, 4.652386, 5.853662, 
    7.579349, 9.558334, 11.55515, 11.73987, 12.24433, 12.31939,
  2.664953, 3.371697, 4.440101, 5.876518, 8.048529, 10.8736, 16.4807, 
    16.11559, 16.05757, 15.88935, 15.49996, 15.4575, 16.41455, 18.60816, 
    21.8139, 25.74877, 30.19903, 27.82057, 27.93264, 27.25346,
  1.958305, 3.50366, 5.977983, 9.282141, 13.83651, 19.33629, 29.32314, 
    29.03934, 29.07602, 28.89136, 28.31006, 28.13081, 29.2514, 31.95641, 
    35.91059, 40.81615, 46.6251, 41.46606, 41.02142, 39.59028,
  -1.727365, 0.8310251, 5.078748, 10.76291, 18.25363, 27.04639, 41.53117, 
    42.58725, 43.47133, 43.586, 42.84328, 42.30365, 43.07615, 45.43468, 
    48.89108, 53.14753, 58.51481, 50.72847, 49.44027, 47.26572,
  -8.954659, -5.291144, 0.9461975, 9.310365, 20.0501, 32.61015, 50.92553, 
    55.32926, 58.45046, 59.53365, 58.75495, 57.49834, 57.07478, 57.71977, 
    58.81231, 60.15406, 62.60285, 53.35073, 50.68176, 47.72026,
  -19.51943, -14.88676, -6.861911, 3.92928, 17.62671, 33.94375, 53.88073, 
    64.27482, 71.91817, 75.23905, 74.68114, 72.03735, 68.95051, 65.8065, 
    62.10393, 57.96612, 54.78806, 47.16319, 42.32716, 38.48795,
  -30.55288, -25.62224, -16.91859, -4.94138, 10.68906, 30.31975, 49.03636, 
    64.59409, 76.57282, 82.57846, 82.96086, 79.50809, 73.87344, 66.55871, 
    57.42559, 47.09581, 37.37708, 34.14541, 25.80407, 20.63282,
  -39.8948, -35.52176, -27.68654, -16.57255, -1.363215, 19.03912, 36.21303, 
    52.38259, 65.41076, 72.87914, 74.63914, 71.75087, 65.23428, 55.53991, 
    43.1028, 29.1264, 15.61026, 12.82065, 1.925284, -4.104444,
  -47.91685, -44.65023, -38.80272, -30.41664, -18.61416, -2.101218, 16.10036, 
    29.5574, 41.10824, 48.29426, 50.39931, 47.70861, 40.75157, 30.29163, 
    17.50934, 3.954396, -8.65477, -19.08495, -28.874, -34.14639,
  -55.22511, -53.26353, -49.83485, -45.02737, -38.34659, -29.16906, 
    -9.008943, -1.761326, 4.89319, 9.115718, 10.01649, 7.350761, 1.368575, 
    -6.968173, -16.35839, -25.63395, -33.72564, -55.54978, -61.77536, -65.2825,
  -62.53136, -61.71577, -60.42729, -58.95439, -57.49697, -56.59324, 
    -35.12228, -35.90551, -36.59852, -37.55915, -39.09142, -41.48574, 
    -44.74864, -48.42105, -51.99606, -55.16397, -57.53818, -90.26324, 
    -92.15633, -93.53811,
  -69.74883, -69.72993, -69.90387, -70.82938, -73.47494, -79.42082, 
    -57.93806, -65.58568, -72.96185, -78.7487, -82.43266, -84.22176, 
    -84.51704, -83.68458, -82.10131, -80.10483, -77.79877, -118.0491, 
    -116.1017, -115.4771,
  -75.76578, -76.21257, -77.16772, -79.40481, -84.48679, -94.50666, 
    -73.95766, -84.82791, -95.23348, -102.9389, -107.2255, -108.5134, 
    -107.5227, -104.8978, -101.1418, -96.68874, -91.9653, -135.3745, 
    -130.8179, -128.6305,
  -78.91267, -79.63683, -80.94291, -83.64637, -89.55829, -100.7131, -81.6423, 
    -91.93498, -101.5724, -108.3939, -111.996, -113.1293, -112.6233, 
    -110.8328, -107.7252, -103.3836, -98.3962, -140.8416, -135.1368, -132.0038,
  -77.79032, -78.71641, -80.17516, -82.80597, -88.28461, -98.24164, -81.3409, 
    -89.10466, -96.18712, -101.0256, -103.5632, -104.707, -105.237, 
    -105.1369, -103.7871, -100.8105, -96.78735, -134.8603, -129.3903, 
    -126.0047,
  -71.89275, -72.93282, -74.37428, -76.5162, -80.61183, -87.83702, -74.22124, 
    -79.89375, -84.80025, -87.95708, -89.57043, -90.50397, -91.43291, 
    -92.23038, -92.09206, -90.38941, -87.5818, -118.7191, -114.7468, -111.8665,
  -61.64122, -62.64447, -63.81977, -65.0298, -66.92556, -70.3405, -61.07608, 
    -66.94012, -71.61501, -74.05221, -74.83157, -74.83986, -74.79147, 
    -74.83215, -74.47487, -73.17902, -71.24721, -93.96004, -92.74217, 
    -91.23203,
  -48.6263, -49.26488, -49.76266, -49.83259, -49.84393, -50.48108, -45.77506, 
    -49.34517, -52.3597, -54.00345, -54.63351, -54.83052, -55.11094, 
    -55.63912, -56.11324, -56.0977, -55.72768, -68.76385, -69.27382, -68.75311,
  -32.78158, -32.92029, -32.68797, -31.89833, -30.87187, -30.19113, -27.9965, 
    -28.15409, -28.80796, -29.56964, -30.35901, -31.36231, -32.76819, 
    -34.52396, -36.31217, -37.76334, -38.88173, -44.82767, -45.55958, -45.3995,
  -13.70377, -13.50742, -12.90668, -11.75581, -10.14503, -8.443991, 
    -6.682826, -5.835516, -5.690591, -6.010222, -6.717126, -7.919562, 
    -9.623322, -11.5973, -13.51622, -15.14572, -16.44324, -18.48131, 
    -19.21223, -19.46359,
  5.855795, 5.739593, 5.387968, 4.785368, 4.104611, 3.542658, 3.825698, 
    3.155673, 2.934653, 2.987202, 3.284466, 4.018037, 5.348554, 7.215276, 
    9.372635, 11.58192, 13.69905, 14.1232, 14.79937, 14.98785,
  13.36187, 13.68183, 13.90033, 13.91653, 14.08323, 14.5514, 17.73631, 
    15.89958, 15.12953, 15.04959, 15.44046, 16.6299, 18.95641, 22.35422, 
    26.41191, 30.8069, 35.42107, 33.72525, 34.21072, 33.78613,
  18.51889, 19.37243, 20.40884, 21.46903, 23.04277, 25.19405, 31.65324, 
    29.43601, 28.49291, 28.34213, 28.7098, 30.11689, 33.08373, 37.50997, 
    42.78233, 48.48428, 54.62295, 50.74521, 50.85861, 49.80118,
  19.87854, 21.40878, 23.60909, 26.27599, 29.97769, 34.70381, 44.71765, 
    43.5962, 43.31095, 43.33378, 43.53853, 44.7429, 47.6804, 52.20054, 
    57.46446, 62.97077, 68.98235, 63.27542, 62.70379, 60.9962,
  16.11338, 18.47042, 22.18721, 27.00225, 33.50219, 41.72776, 55.03945, 
    57.31233, 59.25755, 60.12391, 60.1224, 60.51714, 62.33628, 65.41511, 
    68.74603, 71.84475, 75.35777, 69.06715, 67.23426, 64.80558,
  6.460521, 9.692077, 15.06547, 22.23518, 31.77754, 44.07557, 59.34343, 
    67.96523, 74.74718, 77.87157, 77.77718, 76.38814, 75.31847, 74.64675, 
    73.45692, 71.49079, 69.76059, 65.55745, 61.59363, 58.30383,
  -7.122476, -3.362497, 3.130818, 12.09457, 24.26949, 40.58262, 56.13877, 
    70.76467, 82.59223, 88.66772, 89.25626, 86.54095, 82.42181, 77.21778, 
    70.39788, 62.18013, 53.98354, 53.66079, 46.08971, 41.3777,
  -22.44437, -18.76476, -12.25938, -3.01872, 9.927094, 28.01892, 43.78629, 
    60.17101, 73.99219, 82.11127, 84.19798, 81.72153, 76.02701, 67.52658, 
    56.42074, 43.62558, 30.91572, 30.36727, 19.80522, 13.99333,
  -38.77833, -35.68451, -30.20704, -22.44887, -11.58016, 3.812432, 21.5744, 
    35.87348, 48.82211, 57.22942, 59.91294, 57.35737, 50.43026, 40.04419, 
    27.36016, 13.80649, 1.026303, -7.750523, -17.60755, -22.84733,
  -55.03945, -52.79498, -48.88678, -43.58829, -36.6305, -27.51716, -7.46479, 
    0.3284949, 7.854525, 12.94829, 14.30708, 11.63492, 5.333769, -3.476515, 
    -13.40106, -23.21017, -31.72563, -52.89594, -59.08205, -62.53967,
  -70.19921, -68.77478, -66.37561, -63.52829, -60.75194, -58.88718, 
    -37.10194, -37.67567, -38.3736, -39.37234, -40.91322, -43.3826, -46.924, 
    -51.12196, -55.38316, -59.1764, -61.84853, -95.00439, -96.56904, -97.79725,
  -82.94464, -82.15924, -80.87848, -79.85738, -80.35369, -84.26939, 
    -61.49904, -68.43768, -75.72958, -81.72984, -85.61716, -87.69163, 
    -88.55612, -88.6176, -88.08246, -86.96116, -85.07444, -126.5255, 
    -124.2192, -123.4157,
  -91.79831, -91.49007, -90.95129, -91.03579, -93.47072, -100.6025, 
    -77.56625, -86.89053, -96.49364, -103.9793, -108.4302, -110.3469, 
    -110.4543, -109.2152, -106.8493, -103.4823, -99.37366, -144.3025, 
    -139.6161, -137.3412,
  -95.53635, -95.6254, -95.61967, -96.28569, -99.45085, -107.3466, -84.87334, 
    -93.28976, -101.732, -108.107, -111.9575, -113.9988, -114.8222, 
    -114.4435, -112.5655, -109.1052, -104.6329, -148.5876, -143.0216, 
    -139.9484,
  -93.55219, -93.97942, -94.3787, -95.26097, -98.21319, -105.0447, -84.28994, 
    -90.582, -96.72499, -101.3224, -104.2953, -106.3773, -108.0078, 
    -108.8451, -108.1293, -105.4907, -101.5925, -141.0571, -135.892, -132.7013,
  -85.96571, -86.59959, -87.18816, -87.8954, -89.85158, -94.4082, -76.88407, 
    -81.95084, -86.68554, -90.05206, -92.15777, -93.70541, -95.16677, 
    -96.23641, -96.078, -94.15948, -91.02451, -123.4975, -119.8379, -117.225,
  -73.48742, -74.11964, -74.55705, -74.57935, -74.75142, -76.08646, 
    -63.24706, -69.33281, -74.84768, -77.99997, -79.0498, -78.99788, 
    -78.75919, -78.50735, -77.72284, -75.90623, -73.32726, -97.4886, 
    -96.39326, -95.11646,
  -57.69815, -58.04831, -58.00233, -57.22858, -56.01246, -55.12824, 
    -47.54731, -51.44735, -55.21072, -57.45103, -58.30301, -58.41224, 
    -58.4456, -58.60822, -58.57875, -57.94736, -56.79801, -71.22903, 
    -71.70327, -71.33463,
  -38.64819, -38.62993, -38.11859, -36.8945, -35.16206, -33.45092, -29.24161, 
    -29.32894, -30.06014, -31.07851, -32.24781, -33.55907, -35.0526, 
    -36.63474, -38.03083, -38.95218, -39.42113, -46.30469, -46.99223, 
    -46.91765,
  -16.19345, -15.9391, -15.25225, -13.98118, -12.11821, -9.882509, -7.078318, 
    -5.529467, -4.935811, -5.359741, -6.630142, -8.460152, -10.52767, 
    -12.54186, -14.30298, -15.71543, -16.79266, -19.03098, -19.74169, 
    -20.01045,
  11.12651, 10.83718, 10.12783, 8.9271, 7.31612, 5.467747, 4.190614, 
    2.266345, 1.317763, 1.404925, 2.401477, 4.136312, 6.375374, 8.835114, 
    11.26137, 13.51937, 15.57576, 16.15355, 16.89504, 17.14089,
  25.89302, 25.80096, 25.17995, 23.84805, 22.05586, 20.02875, 20.19798, 
    16.36251, 14.38922, 14.25331, 15.63416, 18.35004, 22.15273, 26.58816, 
    31.13504, 35.53778, 39.82938, 38.73816, 39.3912, 39.13744,
  37.72787, 37.89648, 37.54717, 36.43976, 35.00108, 33.50493, 35.51407, 
    30.66545, 28.09309, 27.76883, 29.35348, 32.75286, 37.73167, 43.64824, 
    49.68542, 55.45742, 61.12427, 58.41739, 58.7633, 57.95831,
  44.79644, 45.31965, 45.50858, 45.12885, 44.79351, 44.87462, 49.14378, 
    44.90734, 42.63937, 42.33175, 43.87517, 47.4356, 52.86649, 59.3451, 
    65.74379, 71.54945, 77.11564, 73.25596, 72.92432, 71.50632,
  45.19948, 46.20808, 47.27939, 48.23211, 49.86381, 52.77319, 59.50225, 
    58.25412, 57.87644, 58.18562, 59.52062, 62.51548, 67.23723, 72.76052, 
    77.73293, 81.60043, 84.96059, 81.10517, 79.50403, 77.37789,
  37.26181, 38.89082, 41.17615, 43.98751, 48.27955, 55.1067, 64.07083, 
    68.67807, 72.65684, 74.88661, 76.02816, 77.40311, 79.60467, 81.91416, 
    83.04874, 82.60503, 81.3995, 79.3596, 75.75145, 72.81318,
  21.66881, 23.89883, 27.45811, 32.30676, 39.51602, 50.52064, 61.518, 
    71.96564, 80.55318, 85.16995, 86.61981, 86.65798, 86.09713, 84.39748, 
    80.62856, 74.81651, 68.19508, 68.55293, 61.79865, 57.57689,
  0.04271889, 2.660983, 7.113199, 13.40199, 22.57612, 36.17237, 49.36931, 
    62.14833, 72.56667, 78.43061, 80.68649, 80.80251, 78.84958, 74.14338, 
    66.39061, 56.3261, 45.73358, 45.23115, 35.76011, 30.48829,
  -25.95173, -23.23117, -18.50307, -11.92712, -2.813111, 10.06841, 26.43958, 
    38.3674, 48.30778, 54.05434, 56.32586, 56.04709, 52.61401, 45.55943, 
    35.51227, 23.86012, 12.46076, 5.020036, -3.965617, -8.741941,
  -52.89085, -50.34403, -45.88395, -39.94978, -32.542, -23.42006, -4.128988, 
    3.274342, 9.423293, 12.82045, 13.78681, 12.52941, 8.233021, 0.9054556, 
    -8.268161, -17.76507, -26.05503, -44.33893, -49.84728, -52.89228,
  -77.08387, -74.92303, -71.10053, -66.31899, -61.37305, -57.30731, 
    -35.55848, -34.29457, -33.75581, -34.06151, -35.23222, -37.72914, 
    -41.96793, -47.47219, -53.22518, -58.19867, -61.48923, -91.10095, 
    -92.07417, -92.93323,
  -95.60562, -93.97049, -90.99446, -87.52327, -84.98239, -85.39599, 
    -61.53647, -65.03756, -68.95012, -72.21174, -75.16749, -78.66366, 
    -82.44225, -85.69495, -87.85174, -88.54803, -87.61015, -125.8752, 
    -123.1544, -122.0884,
  -106.9161, -105.8774, -103.8369, -101.6187, -100.9554, -104.2447, -78.894, 
    -84.31635, -89.8045, -94.02745, -97.73361, -101.7953, -105.4025, 
    -107.4796, -107.6016, -105.7875, -102.4926, -145.0194, -140.2101, 
    -137.8466,
  -110.7312, -110.2824, -109.1519, -107.9935, -108.4994, -112.9066, 
    -87.22113, -92.30766, -97.09164, -100.7711, -104.3962, -108.5928, 
    -112.2943, -114.2479, -113.8578, -111.1876, -107.0749, -149.3734, 
    -143.9622, -140.9885,
  -107.502, -107.5389, -107.1439, -106.7061, -107.6152, -111.6732, -87.29993, 
    -91.45013, -95.04681, -97.88564, -101.0085, -104.7485, -108.1501, 
    -110.0485, -109.6914, -107.0125, -102.9126, -141.3533, -136.4919, 
    -133.5446,
  -98.01415, -98.32743, -98.32131, -98.09299, -98.60624, -101.2207, 
    -80.10278, -84.26228, -87.7788, -90.31227, -92.62198, -95.02029, 
    -97.11119, -98.18779, -97.55807, -95.00167, -91.18594, -123.2588, 
    -119.8371, -117.5099,
  -83.26402, -83.57918, -83.49062, -82.80865, -82.05726, -82.32458, 
    -66.33459, -72.15332, -77.56608, -80.69067, -81.78443, -81.70155, 
    -81.16766, -80.29472, -78.67024, -75.97855, -72.42263, -96.93981, 
    -95.72493, -94.6142,
  -64.89059, -64.98791, -64.56137, -63.34994, -61.62987, -60.19062, -50.081, 
    -54.00474, -57.82645, -60.05186, -60.81459, -60.70438, -60.3231, 
    -59.84675, -58.99519, -57.45784, -55.22345, -70.5493, -70.69444, -70.3722,
  -43.14316, -42.98294, -42.28541, -40.88552, -38.9352, -36.85473, -30.92078, 
    -31.05733, -31.56346, -32.34485, -33.48645, -34.83645, -36.20836, 
    -37.41441, -38.21357, -38.40132, -37.98283, -45.64414, -46.08117, 
    -46.00901,
  -18.10965, -17.77335, -16.98455, -15.64882, -13.73872, -11.34596, 
    -7.852421, -5.827647, -4.692091, -4.924373, -6.444824, -8.648508, 
    -10.90845, -12.87339, -14.42918, -15.56867, -16.32937, -18.68265, 
    -19.25728, -19.48216,
  13.42813, 13.04794, 12.17689, 10.75331, 8.834326, 6.555789, 4.667517, 
    2.211428, 0.8663781, 0.8723874, 2.101475, 4.205895, 6.758179, 9.380908, 
    11.82411, 13.99444, 15.89956, 16.46578, 17.14705, 17.37068,
  31.29523, 31.02575, 30.08359, 28.29323, 25.86374, 23.00066, 21.9292, 
    17.28554, 14.63944, 14.25481, 15.87037, 19.08231, 23.34144, 27.9988, 
    32.48651, 36.58421, 40.39217, 39.44756, 39.99112, 39.72844,
  45.90022, 45.80231, 44.95508, 43.11439, 40.65789, 37.87812, 37.97202, 
    32.02415, 28.52154, 27.81862, 29.68826, 33.75752, 39.37275, 45.59812, 
    51.53083, 56.82487, 61.72155, 59.3376, 59.49889, 58.681,
  55.24754, 55.4025, 54.88231, 53.43856, 51.64492, 49.9517, 51.6149, 
    45.90868, 42.42127, 41.61758, 43.55281, 48.04372, 54.38111, 61.33788, 
    67.67185, 72.9264, 77.53165, 74.13836, 73.51415, 72.05685,
  57.31069, 57.8281, 57.93732, 57.44711, 57.14902, 57.78056, 61.34901, 
    58.03914, 55.97144, 55.58604, 57.46143, 61.78128, 67.84473, 74.18641, 
    79.31982, 82.77235, 85.19849, 81.74282, 79.77425, 77.58913,
  50.22804, 51.235, 52.30121, 53.3153, 55.27534, 59.38823, 65.17919, 
    66.73639, 68.12891, 69.22659, 71.08994, 74.40292, 78.64791, 82.38823, 
    84.20911, 83.83419, 82.15515, 79.70535, 75.88761, 72.959,
  34.29094, 35.85404, 38.10101, 41.00784, 45.65446, 53.49096, 61.9716, 
    68.37169, 73.24537, 75.89655, 77.92985, 80.43893, 82.76895, 83.40732, 
    81.23066, 76.42175, 70.37145, 69.01266, 62.67192, 58.70004,
  10.81198, 12.87512, 16.22927, 20.85918, 27.7148, 38.1023, 49.41028, 
    57.79168, 63.65415, 66.45042, 68.57146, 71.21729, 72.84308, 71.44923, 
    66.31911, 58.28886, 49.39611, 47.1881, 38.77976, 33.99595,
  -18.38668, -15.97593, -11.85155, -6.197721, 1.540891, 12.27322, 27.16221, 
    35.539, 41.14043, 43.43611, 45.01014, 46.93565, 47.10832, 43.57089, 
    36.34537, 26.86462, 17.25733, 10.12199, 2.244426, -2.014499,
  -49.11974, -46.58903, -42.13445, -36.20325, -28.88284, -20.09824, 
    -1.814556, 4.460468, 8.515539, 9.908045, 10.39612, 10.47928, 8.398238, 
    3.114124, -4.570481, -13.01228, -20.50965, -35.91563, -40.72154, -43.37224,
  -76.67981, -74.32523, -70.07256, -64.59547, -58.68138, -53.3018, -32.02391, 
    -29.06765, -27.31296, -26.9225, -27.69356, -30.02348, -34.46264, 
    -40.52917, -46.94973, -52.43703, -56.09211, -81.04333, -81.74383, 
    -82.37448,
  -97.46993, -95.57663, -92.0332, -87.61877, -83.66486, -81.98838, -58.17137, 
    -58.39948, -58.82812, -59.34346, -61.25367, -65.6364, -71.57172, 
    -77.2273, -81.32383, -83.29447, -83.16055, -116.297, -113.5272, -112.3636,
  -109.8701, -108.615, -106.1027, -103.0767, -101.1251, -102.4304, -76.81863, 
    -78.99303, -80.58633, -81.58687, -84.24538, -89.71547, -96.00249, 
    -100.6294, -102.5403, -101.7724, -99.06347, -136.9963, -132.2224, 
    -129.8529,
  -113.8946, -113.3009, -111.8749, -110.2055, -109.8299, -112.814, -86.63421, 
    -89.39155, -91.02482, -92.01595, -94.89136, -100.4054, -106.1981, 
    -109.8284, -110.4004, -108.1712, -104.2254, -142.8835, -137.5586, 
    -134.6524,
  -110.352, -110.2959, -109.7517, -109.0826, -109.5485, -112.8264, -87.79552, 
    -90.66922, -92.14265, -93.053, -95.66048, -100.2761, -104.8518, 
    -107.4412, -107.2589, -104.4924, -100.1981, -135.9912, -131.233, -128.4042,
  -100.2884, -100.5306, -100.4584, -100.195, -100.6334, -103.0492, -81.19279, 
    -84.7775, -87.0107, -88.27802, -90.20794, -93.0087, -95.51574, -96.59552, 
    -95.64753, -92.68472, -88.42787, -118.777, -115.371, -113.1565,
  -84.86576, -85.10372, -84.96742, -84.3568, -83.83597, -84.48306, -67.7658, 
    -73.05775, -77.55807, -79.94211, -80.86707, -80.93959, -80.39921, 
    -79.19408, -77.04861, -73.82829, -69.68323, -93.37018, -91.90781, 
    -90.80401,
  -65.83545, -65.87507, -65.43613, -64.35713, -62.97847, -62.07711, 
    -51.27878, -54.93859, -58.15947, -59.84215, -60.38672, -60.24033, 
    -59.71894, -58.89005, -57.5409, -55.46891, -52.59964, -67.82915, 
    -67.61657, -67.23276,
  -43.5924, -43.40527, -42.72361, -41.44796, -39.75322, -38.01208, -31.65928, 
    -31.93623, -32.17658, -32.49403, -33.28372, -34.45192, -35.675, 
    -36.64628, -37.1029, -36.8765, -35.94885, -43.77246, -43.96217, -43.83509,
  -18.29669, -17.92945, -17.11201, -15.79475, -13.98504, -11.77207, 
    -8.309644, -6.414628, -5.165468, -5.09456, -6.316972, -8.353409, 
    -10.55023, -12.46995, -13.94355, -14.95239, -15.53101, -17.87289, 
    -18.32335, -18.49658,
  14.63267, 14.19594, 13.23512, 11.71337, 9.694975, 7.304052, 5.203221, 
    2.580209, 1.018777, 0.8586901, 2.034292, 4.172362, 6.772101, 9.394476, 
    11.76336, 13.78515, 15.4833, 15.97141, 16.53847, 16.70885,
  34.08175, 33.71881, 32.6342, 30.68483, 28.07211, 24.98692, 23.36368, 
    18.4784, 15.41253, 14.63674, 16.05267, 19.23936, 23.5072, 28.06491, 
    32.27407, 35.90591, 39.09288, 38.12373, 38.42845, 38.08426,
  50.02228, 49.79748, 48.74813, 46.65574, 43.87175, 40.67965, 39.80181, 
    33.44512, 29.29612, 28.01913, 29.62878, 33.71091, 39.37597, 45.45808, 
    50.9509, 55.50626, 59.40754, 57.03518, 56.80969, 55.86834,
  60.36768, 60.36111, 59.56062, 57.72066, 55.3646, 52.94137, 53.11621, 
    46.60703, 42.12011, 40.56308, 42.29994, 47.0285, 53.63974, 60.55558, 
    66.40665, 70.76297, 74.10384, 70.66679, 69.49654, 67.86523,
  63.0979, 63.40756, 63.1228, 62.02333, 60.82344, 60.24885, 61.81808, 
    56.89387, 53.15617, 51.72005, 53.56514, 58.61396, 65.48532, 72.17014, 
    77.02855, 79.67062, 80.82767, 76.97955, 74.39752, 72.02487,
  56.45289, 57.18288, 57.69633, 57.83036, 58.48565, 60.78955, 64.44808, 
    62.99139, 61.48166, 60.92941, 62.99883, 67.88376, 73.91246, 78.7959, 
    80.93849, 80.25476, 77.82054, 73.82815, 69.6626, 66.66782,
  40.77686, 42.00269, 43.55371, 45.31949, 48.21767, 53.45649, 60.08616, 
    62.00108, 62.52539, 62.58603, 64.73872, 69.53905, 74.77945, 77.72588, 
    76.95203, 72.89812, 67.27071, 63.05214, 57.16659, 53.45825,
  17.37421, 19.08405, 21.70572, 25.12055, 30.04673, 37.36786, 46.90401, 
    50.19448, 50.91574, 50.29295, 51.93832, 56.82285, 61.97308, 63.96379, 
    61.48749, 55.50964, 48.40831, 43.74314, 36.6095, 32.40607,
  -11.99664, -9.896881, -6.384953, -1.690532, 4.562081, 12.86562, 25.97461, 
    30.11465, 31.13887, 30.1844, 31.02438, 34.73436, 38.22475, 38.25374, 
    34.08111, 27.08118, 19.61687, 12.48322, 5.950211, 2.295833,
  -43.24358, -40.91838, -36.82053, -31.35296, -24.63302, -16.74136, 
    0.02973527, 4.59485, 6.409999, 6.101265, 6.263091, 7.500843, 7.577695, 
    4.654291, -1.014508, -7.87737, -14.19111, -26.43868, -30.49271, -32.74794,
  -71.64943, -69.37997, -65.21635, -59.71488, -53.52974, -47.44539, 
    -27.29445, -23.04942, -20.43318, -19.51682, -19.81248, -21.60891, 
    -25.58309, -31.41452, -37.79069, -43.31326, -47.17003, -66.41364, 
    -67.03127, -67.5208,
  -93.43726, -91.54973, -87.94083, -83.24648, -78.56666, -75.33038, 
    -52.45988, -49.53676, -46.79741, -44.95026, -45.69908, -50.16066, 
    -57.23796, -64.54655, -70.16566, -73.2614, -74.03036, -100.2691, 
    -97.71999, -96.56972,
  -106.7392, -105.467, -102.8759, -99.58839, -96.9474, -96.74387, -72.0974, 
    -70.98807, -68.75601, -66.6536, -67.90213, -73.90864, -82.15601, 
    -89.07887, -92.79871, -93.19363, -91.24111, -122.4887, -117.9251, 
    -115.6208,
  -111.4074, -110.8083, -109.3727, -107.6187, -106.8801, -108.9269, 
    -83.69667, -84.12286, -82.55053, -80.68319, -82.26139, -88.39264, 
    -95.96071, -101.3587, -103.1048, -101.5, -97.84538, -130.9215, -125.7203, 
    -122.8954,
  -108.2323, -108.1889, -107.717, -107.166, -107.6568, -110.6634, -86.41263, 
    -88.02094, -87.2673, -85.94913, -87.49129, -92.51131, -98.18751, 
    -101.6655, -101.8904, -99.20994, -94.81116, -126.4151, -121.704, -118.9636,
  -98.3477, -98.6129, -98.66995, -98.68502, -99.49068, -102.2232, -80.8539, 
    -83.74018, -84.44411, -84.09619, -85.26043, -88.28142, -91.30811, 
    -92.616, -91.55659, -88.33862, -83.72406, -111.2282, -107.7376, -105.5789,
  -83.04288, -83.29691, -83.3035, -83.07023, -83.22272, -84.77694, -68.15946, 
    -72.58356, -75.65762, -76.89586, -77.54405, -77.9758, -77.74876, 
    -76.46699, -73.96339, -70.32181, -65.66001, -87.72141, -85.8956, -84.72795,
  -64.20633, -64.2672, -63.97314, -63.27447, -62.59743, -62.67496, -51.67944, 
    -54.79475, -57.02826, -57.90185, -58.20729, -58.21885, -57.80434, 
    -56.8057, -55.07443, -52.55339, -49.12569, -63.76126, -63.10188, -62.59839,
  -42.37735, -42.21383, -41.64386, -40.63638, -39.4065, -38.28633, -31.87549, 
    -32.26788, -32.19064, -31.95284, -32.27705, -33.20407, -34.29738, 
    -35.09553, -35.2816, -34.71478, -33.35151, -41.09328, -40.99403, -40.78218,
  -17.74357, -17.3694, -16.56383, -15.31855, -13.69228, -11.81156, -8.643315, 
    -7.128163, -5.96411, -5.570166, -6.25236, -7.844142, -9.821644, 
    -11.66631, -13.0874, -14.00592, -14.43675, -16.72418, -17.04516, -17.1619,
  14.75161, 14.29697, 13.32061, 11.81485, 9.871311, 7.629689, 5.663554, 
    3.217464, 1.644393, 1.2738, 2.137335, 3.985664, 6.376313, 8.846911, 
    11.06676, 12.90213, 14.36742, 14.73976, 15.16585, 15.26779,
  34.27055, 33.89924, 32.84061, 30.99158, 28.56638, 25.75367, 24.165, 
    19.53834, 16.32689, 15.09026, 15.94575, 18.64122, 22.51803, 26.70688, 
    30.47633, 33.54296, 36.03419, 34.90731, 34.88747, 34.41279,
  50.15015, 49.92857, 48.93797, 46.99457, 44.43669, 41.52717, 40.47441, 
    34.29716, 29.78854, 27.81212, 28.70077, 32.21855, 37.43719, 43.03534, 
    47.87716, 51.55714, 54.35524, 51.74994, 51.00694, 49.86861,
  60.28134, 60.2915, 59.56844, 57.8728, 55.67046, 53.3574, 53.00637, 
    46.26593, 40.99364, 38.45813, 39.4385, 43.76023, 50.11924, 56.6489, 
    61.80921, 65.1322, 67.1052, 63.23734, 61.38298, 59.50051,
  62.78373, 63.11562, 62.89314, 61.85188, 60.58329, 59.69212, 60.3154, 
    54.21665, 48.87749, 46.03465, 47.19673, 52.3021, 59.49839, 66.25745, 
    70.70187, 72.45347, 72.30758, 67.50192, 64.23198, 61.62554,
  56.2378, 56.96448, 57.45698, 57.45531, 57.66883, 58.97153, 61.53094, 
    57.30571, 52.8425, 50.19246, 51.71872, 57.46643, 64.87291, 70.76418, 
    73.20184, 72.21751, 69.10446, 62.86954, 58.40673, 55.36008,
  41.39396, 42.55109, 43.91531, 45.21995, 47.10544, 50.3632, 55.9514, 
    53.51454, 49.74684, 46.9578, 48.51082, 54.75907, 62.39561, 67.5079, 
    68.15118, 64.91174, 59.82792, 52.24677, 46.95523, 43.57327,
  19.79812, 21.33797, 23.56166, 26.17768, 29.58431, 34.15861, 42.35495, 
    40.80059, 36.94349, 33.32417, 34.14633, 40.25946, 47.97709, 52.84904, 
    52.86808, 48.94356, 43.68747, 36.37018, 30.64443, 27.08831,
  -6.999138, -5.179044, -2.239161, 1.504554, 6.211411, 11.9553, 23.28333, 
    23.41139, 20.75326, 17.51038, 17.72065, 22.34408, 28.04748, 30.94636, 
    29.5816, 25.0578, 19.79756, 12.50371, 7.387288, 4.361373,
  -35.67554, -33.68583, -30.20786, -25.59784, -19.98819, -13.59944, 1.177412, 
    3.739887, 3.67249, 2.302505, 2.378328, 4.452964, 6.255728, 5.5699, 
    2.089835, -2.941539, -7.873024, -17.05013, -20.384, -22.2889,
  -62.40727, -60.44573, -56.80551, -51.8904, -46.16887, -40.22185, -22.11946, 
    -17.4999, -14.68989, -13.51015, -13.23888, -14.08905, -16.85757, 
    -21.53979, -27.06703, -32.11105, -35.95192, -49.16612, -49.88518, 
    -50.34369,
  -83.80297, -82.14448, -78.90104, -74.51856, -69.79294, -65.71287, 
    -44.99369, -39.90224, -35.17932, -31.82075, -31.37113, -34.87986, 
    -41.53646, -49.11441, -55.42525, -59.32709, -61.03062, -79.3616, 
    -77.33031, -76.33121,
  -97.72462, -96.60701, -94.26582, -91.15995, -88.31493, -87.03716, 
    -64.72124, -60.88442, -55.74376, -51.26731, -50.88404, -56.17331, 
    -64.8997, -73.22236, -78.51762, -80.19673, -79.26186, -102.2248, 
    -98.13419, -96.00412,
  -103.4798, -102.9939, -101.7731, -100.2324, -99.4465, -100.7921, -77.94038, 
    -76.16427, -71.79638, -67.36842, -67.23792, -72.95742, -81.47235, 
    -88.48298, -91.67558, -91.04283, -87.96249, -113.6964, -108.7438, 
    -106.0472,
  -101.4484, -101.5055, -101.2685, -101.0501, -101.7962, -104.6991, 
    -82.55826, -82.77305, -79.8516, -76.31009, -76.38125, -81.19757, 
    -87.73972, -92.35509, -93.39943, -91.1436, -86.84751, -112.7374, 
    -108.068, -105.4052,
  -92.61228, -92.97753, -93.30491, -93.78563, -95.16856, -98.38535, 
    -78.54501, -80.43581, -79.44642, -77.36502, -77.51553, -80.56597, 
    -84.24724, -86.15223, -85.34611, -82.12646, -77.29211, -100.8113, 
    -97.15603, -95.00597,
  -78.28181, -78.62923, -78.92199, -79.26294, -80.32056, -82.96999, 
    -67.02619, -70.18594, -71.50179, -71.38728, -71.6836, -72.65147, 
    -73.14354, -72.20317, -69.62978, -65.72829, -60.63147, -80.26343, 
    -77.96613, -76.67134,
  -60.46043, -60.60839, -60.58095, -60.43076, -60.6556, -61.88514, -50.93543, 
    -53.1867, -54.18161, -54.12689, -54.21831, -54.59965, -54.62201, 
    -53.75206, -51.8344, -48.97794, -45.06289, -58.61775, -57.42615, -56.75112,
  -39.8229, -39.72588, -39.34536, -38.71109, -38.07262, -37.7067, -31.40704, 
    -31.78072, -31.33264, -30.55838, -30.44128, -31.16166, -32.19704, 
    -32.91782, -32.92649, -32.10074, -30.37205, -37.80433, -37.38039, 
    -37.05941,
  -16.5914, -16.23132, -15.47613, -14.35752, -12.99083, -11.54757, -8.814144, 
    -7.764699, -6.789397, -6.14407, -6.242836, -7.238595, -8.848494, 
    -10.55164, -11.92595, -12.79172, -13.11726, -15.32176, -15.51995, 
    -15.58243,
  13.07461, 12.66023, 11.7906, 10.50234, 8.93906, 7.274103, 5.935304, 
    4.14535, 2.81802, 2.149811, 2.296903, 3.307284, 4.995319, 6.973969, 
    8.841766, 10.36123, 11.48474, 11.66876, 11.88378, 11.88248,
  30.09473, 29.85243, 29.10192, 27.78748, 26.13658, 24.31793, 23.44646, 
    19.70617, 16.59189, 14.66744, 14.3567, 15.79928, 18.58844, 21.87708, 
    24.81334, 26.97918, 28.42745, 26.91646, 26.34886, 25.64038,
  43.51387, 43.50404, 42.99471, 41.83102, 40.30885, 38.61176, 38.1997, 
    32.83643, 28.07737, 24.95708, 24.29773, 26.32296, 30.29649, 34.81424, 
    38.54586, 40.91986, 42.12554, 38.89568, 37.30602, 35.82539,
  51.40813, 51.70128, 51.58641, 50.80306, 49.69086, 48.48299, 48.49694, 
    41.9557, 35.71781, 31.44551, 30.58825, 33.45731, 38.79492, 44.46103, 
    48.60233, 50.55692, 50.72443, 45.81523, 42.9575, 40.69449,
  52.38805, 53.0423, 53.46906, 53.30257, 52.89672, 52.5559, 53.19587, 
    45.93207, 38.42649, 33.07687, 32.19786, 36.19489, 43.0571, 49.7065, 
    53.76511, 54.63455, 53.08644, 46.36293, 42.28925, 39.42124,
  45.87037, 46.88669, 47.91877, 48.52398, 49.06822, 49.90794, 52.47914, 
    44.94802, 36.66888, 30.62927, 30.01596, 35.27008, 43.47147, 50.56504, 
    53.84429, 53.10847, 49.77715, 39.86874, 35.34081, 32.37842,
  33.47745, 34.78604, 36.36415, 37.67979, 38.93525, 40.25912, 45.94275, 
    38.42491, 29.74805, 23.20794, 22.66584, 28.71173, 37.81255, 45.22703, 
    48.09056, 46.64095, 43.01733, 30.6715, 26.56323, 23.80777,
  17.1313, 18.58608, 20.53032, 22.38345, 24.0965, 25.44614, 33.06476, 
    26.34159, 18.15017, 11.65236, 10.8519, 16.54729, 25.30827, 32.52073, 
    35.47291, 34.51844, 32.05421, 21.24453, 17.6674, 15.12101,
  -2.182395, -0.7246933, 1.430368, 3.787596, 6.216106, 8.389398, 17.77214, 
    13.64698, 7.91693, 3.088757, 2.587044, 7.104704, 13.76389, 18.90327, 
    20.57221, 19.24874, 16.98655, 9.40449, 6.295326, 4.164265,
  -22.81894, -21.41039, -19.06908, -16.14912, -12.82519, -9.442078, 1.845713, 
    1.530869, -0.4174386, -2.397288, -2.107369, 0.7699621, 4.22969, 6.078385, 
    5.479939, 3.08322, 0.2219431, -4.94559, -7.304948, -8.781443,
  -43.08338, -41.77728, -39.34618, -36.02043, -32.06198, -27.87825, 
    -14.65889, -11.3299, -9.356778, -8.134748, -6.857289, -5.776755, 
    -5.870576, -7.691804, -10.87354, -14.48721, -17.89665, -22.619, 
    -23.67598, -24.24947,
  -61.04253, -59.9677, -57.75671, -54.57916, -50.83639, -47.06813, -32.19227, 
    -26.64372, -21.51445, -17.34745, -15.12915, -15.82599, -19.36509, 
    -24.61716, -29.97689, -34.15891, -37.07331, -43.28713, -42.49103, 
    -41.97082,
  -74.67612, -74.00389, -72.43509, -70.13696, -67.65434, -65.67632, 
    -49.63865, -43.8956, -36.99851, -30.71708, -27.88183, -30.14823, 
    -36.45154, -44.06725, -50.2982, -53.7159, -54.76518, -63.78121, 
    -61.03482, -59.44912,
  -82.3591, -82.19974, -81.56377, -80.62862, -80.01302, -80.47034, -63.78649, 
    -59.52969, -52.54712, -45.53102, -42.65409, -45.91988, -53.44872, 
    -61.42509, -66.69399, -68.15585, -66.72895, -78.93875, -74.85706, 
    -72.55383,
  -83.30766, -83.62743, -83.90808, -84.31251, -85.42953, -87.92419, 
    -71.18464, -69.05885, -63.38803, -57.10489, -54.73851, -58.11059, 
    -64.91631, -71.20408, -74.22777, -73.48164, -70.01508, -84.6266, 
    -80.21524, -77.73343,
  -77.69524, -78.30393, -79.16593, -80.41835, -82.58784, -86.17918, 
    -70.28111, -69.96049, -66.33232, -61.83495, -60.33557, -63.05729, 
    -67.76994, -71.27887, -71.77374, -69.26583, -64.5265, -79.79855, 
    -75.84283, -73.6589,
  -66.47002, -67.05473, -67.92297, -69.24133, -71.63192, -75.59025, 
    -61.45547, -62.00875, -60.42886, -58.22773, -57.87768, -59.75826, 
    -62.02018, -62.62529, -60.81526, -57.02283, -51.49146, -65.81714, 
    -62.62342, -61.03107,
  -51.63659, -52.00092, -52.50907, -53.30723, -54.90923, -57.65992, 
    -46.97461, -47.37823, -46.30508, -44.84089, -44.6441, -45.84491, 
    -47.16085, -47.26751, -45.67891, -42.65644, -38.15601, -49.10946, 
    -46.94001, -45.90879,
  -34.04159, -34.10101, -34.09779, -34.11903, -34.42049, -35.14916, 
    -29.06163, -29.03077, -27.9099, -26.46701, -25.89909, -26.51539, 
    -27.69973, -28.57635, -28.57114, -27.54742, -25.39519, -31.92435, 
    -30.93797, -30.40849,
  -13.98805, -13.68148, -13.06861, -12.24251, -11.39055, -10.70574, 
    -8.671804, -8.197795, -7.489902, -6.661416, -6.128692, -6.273018, 
    -7.162958, -8.475492, -9.720776, -10.54958, -10.79511, -12.82886, 
    -12.86533, -12.85737,
  10.89048, 10.54312, 9.823922, 8.795928, 7.625705, 6.481859, 5.672259, 
    4.369325, 3.248518, 2.429001, 2.108522, 2.484037, 3.556754, 5.062624, 
    6.611955, 7.906958, 8.833337, 8.909674, 9.011368, 8.95602,
  24.78187, 24.6988, 24.28616, 23.49799, 22.53989, 21.52801, 21.26187, 
    18.11171, 15.07754, 12.72899, 11.64757, 12.19174, 14.14356, 16.74162, 
    19.10662, 20.73235, 21.587, 19.80075, 18.901, 18.05064,
  35.29094, 35.51812, 35.49873, 35.06314, 34.43764, 33.70633, 33.90524, 
    29.05567, 24.12358, 20.23927, 18.49894, 19.41764, 22.44334, 26.20371, 
    29.28015, 30.96889, 31.34625, 27.66709, 25.60037, 23.92984,
  40.80137, 41.38273, 41.84812, 41.88873, 41.72464, 41.43856, 42.02298, 
    35.64806, 28.82061, 23.37262, 21.11728, 22.73301, 27.15473, 32.21352, 
    35.87867, 37.28833, 36.69758, 31.0804, 27.76291, 25.3393,
  40.4388, 41.3863, 42.38654, 42.98945, 43.38474, 43.65935, 44.8977, 
    37.14547, 28.51569, 21.58228, 19.01672, 21.65022, 27.73021, 34.13376, 
    38.20064, 39.03481, 37.23257, 29.29771, 25.03442, 22.14224,
  34.24853, 35.49775, 36.97072, 38.11922, 39.1245, 40.03239, 43.45847, 
    34.52151, 24.5637, 16.65506, 14.1747, 17.99701, 25.6074, 32.9757, 
    37.00617, 37.06966, 34.3574, 22.37534, 18.11853, 15.34816,
  24.30655, 25.71589, 27.45628, 28.8733, 29.99017, 30.63731, 37.39187, 
    27.95893, 17.54206, 9.338215, 7.073498, 11.62603, 20.04181, 27.87704, 
    31.97282, 32.04846, 29.86349, 15.08697, 11.8649, 9.574089,
  12.53107, 13.91412, 15.66568, 17.08156, 17.97297, 17.96223, 26.26488, 
    17.91325, 8.600821, 1.217515, -0.6884055, 3.697965, 11.54191, 18.82194, 
    22.85854, 23.57705, 22.85509, 10.33872, 8.072909, 6.159781,
  -0.6011896, 0.6189033, 2.260496, 3.741505, 4.856424, 5.235639, 14.07055, 
    8.504477, 2.044804, -3.070691, -3.954992, -0.06872034, 6.132284, 
    11.50433, 14.21178, 14.43492, 13.79103, 6.096478, 4.15003, 2.548409,
  -14.4733, -13.43036, -11.83416, -10.07105, -8.33103, -6.95313, 2.065724, 
    0.2062765, -2.517587, -4.585881, -4.082031, -0.8736366, 3.18651, 
    6.060103, 6.811485, 5.815422, 4.163379, 1.174703, -0.5911725, -1.824029,
  -28.72004, -27.84012, -26.24269, -24.1263, -21.71178, -19.37987, -10.18849, 
    -8.502677, -7.505885, -6.393353, -4.450748, -2.051411, -0.3111248, 
    -0.09845114, -1.507238, -3.950871, -6.841774, -6.71331, -7.973095, 
    -8.661776,
  -42.62302, -41.9565, -40.51093, -38.35569, -35.7755, -33.22359, -23.6677, 
    -19.40543, -15.18718, -11.0837, -7.825087, -6.39735, -7.163145, 
    -9.782663, -13.41607, -17.06871, -20.44222, -19.27424, -19.42421, 
    -19.32926,
  -54.76816, -54.43067, -53.4606, -51.8696, -49.99803, -48.3349, -38.16586, 
    -32.78737, -26.24589, -19.71972, -15.51742, -15.26311, -18.6122, 
    -23.96326, -29.37231, -33.3264, -35.72829, -35.53445, -34.06979, -33.04145,
  -63.29817, -63.38982, -63.18718, -62.6916, -62.25947, -62.34212, -51.37323, 
    -46.40984, -38.92914, -31.15702, -26.7288, -27.69438, -33.05268, 
    -40.05256, -45.82981, -48.69145, -48.86243, -51.2634, -48.24159, -46.40751,
  -66.61992, -67.13403, -67.75527, -68.48929, -69.66522, -71.61573, -59.8469, 
    -56.28228, -49.40045, -41.9511, -38.14902, -40.00864, -45.98318, 
    -52.67912, -57.04677, -57.81087, -55.50553, -61.1742, -57.26026, -55.02643,
  -64.03324, -64.81639, -66.0091, -67.63859, -70.02756, -73.37059, -61.14308, 
    -59.03121, -53.7981, -48.0077, -45.48496, -47.70912, -52.82797, 
    -57.56544, -59.48992, -58.06055, -53.83389, -62.09927, -58.03507, 
    -55.85148,
  -55.88545, -56.64857, -57.89435, -59.75504, -62.73235, -67.00109, 
    -54.67142, -53.18642, -49.72081, -46.2269, -45.35749, -47.69987, 
    -51.32683, -53.60281, -53.06135, -49.8762, -44.32296, -53.88913, 
    -50.01199, -48.16808,
  -43.95726, -44.48861, -45.36389, -46.73035, -49.03601, -52.38813, -42.0745, 
    -41.00633, -38.55014, -36.19379, -35.772, -37.5272, -39.99081, -41.31403, 
    -40.52438, -37.76661, -33.03907, -41.53262, -38.58387, -37.24723,
  -29.12822, -29.31091, -29.57783, -30.0205, -30.86088, -32.14606, -26.18926, 
    -25.65811, -24.02281, -22.21556, -21.48634, -22.18355, -23.65064, 
    -24.86318, -25.08177, -24.0989, -21.75767, -27.36404, -25.9416, -25.23975,
  -11.77358, -11.52494, -11.05346, -10.48802, -10.03586, -9.853298, 
    -8.222197, -7.964437, -7.352492, -6.499176, -5.775805, -5.544526, 
    -5.976689, -6.931202, -8.006773, -8.796965, -9.018713, -10.89779, 
    -10.83889, -10.79142,
  8.036471, 7.782848, 7.265956, 6.566756, 5.850638, 5.244772, 4.926128, 
    4.019944, 3.054676, 2.118263, 1.42458, 1.239651, 1.694961, 2.669449, 
    3.847812, 4.91256, 5.680148, 5.682305, 5.713202, 5.627731,
  17.89234, 18.00329, 17.98363, 17.77145, 17.51587, 17.24784, 17.49584, 
    14.75614, 11.70603, 8.954595, 7.202949, 6.952757, 8.128317, 10.07436, 
    11.93491, 13.14208, 13.56399, 11.55608, 10.41426, 9.46749,
  24.80552, 25.30005, 25.80987, 26.11835, 26.34882, 26.46382, 27.19025, 
    22.65358, 17.47195, 12.86572, 10.13587, 10.02073, 12.14457, 15.22303, 
    17.80842, 19.0747, 18.94732, 14.91672, 12.5501, 10.77535,
  27.61124, 28.48808, 29.53043, 30.35921, 31.06282, 31.57299, 32.76196, 
    26.46969, 19.1311, 12.6536, 9.078344, 9.388547, 12.78513, 17.22457, 
    20.60485, 21.85739, 21.0148, 14.85594, 11.36866, 8.918692,
  26.01951, 27.22849, 28.73601, 30.01591, 31.12577, 31.9709, 34.069, 
    26.05448, 16.70806, 8.552948, 4.390377, 5.410114, 10.29274, 16.1803, 
    20.3396, 21.56391, 20.12496, 11.26003, 7.14915, 4.383872,
  20.6003, 22.01268, 23.80733, 25.38131, 26.81651, 27.93417, 32.65005, 
    23.00815, 12.208, 3.052671, -1.173364, 0.7620821, 6.995436, 13.99226, 
    18.62234, 19.81619, 18.2712, 4.788365, 0.9921017, -1.505908,
  13.61715, 15.03959, 16.8099, 18.245, 19.33014, 19.74446, 28.08905, 
    17.88457, 6.850708, -2.271641, -6.09343, -3.497078, 3.316759, 10.63621, 
    15.44602, 17.02061, 16.46937, 0.02961588, -2.356207, -4.203173,
  6.735422, 7.977234, 9.449224, 10.43605, 10.7755, 10.09896, 19.67851, 
    10.88547, 1.423848, -6.291145, -9.162306, -6.336373, -0.04164791, 
    6.451399, 10.81708, 12.7504, 13.52231, -0.1654882, -1.306953, -2.660127,
  -0.09702058, 0.8670411, 1.995193, 2.702188, 2.833086, 2.089154, 10.88003, 
    4.724436, -1.883769, -7.036179, -8.276178, -5.165569, 0.1991439, 
    5.184184, 8.244539, 9.46806, 10.06687, 2.359175, 1.402835, 0.2661107,
  -7.043516, -6.330478, -5.406382, -4.671283, -4.285388, -4.533332, 2.489263, 
    -0.5422462, -3.82301, -5.939732, -5.292359, -1.912414, 2.441743, 
    5.877135, 7.481797, 7.512248, 6.868305, 5.690774, 4.491265, 3.490445,
  -14.73655, -14.21795, -13.36076, -12.38568, -11.5154, -11.11787, -6.016884, 
    -6.09536, -6.142767, -5.224718, -2.761251, 0.7255502, 3.982442, 5.909348, 
    6.078585, 4.786854, 2.554827, 6.798625, 5.454484, 4.678567,
  -23.56949, -23.24883, -22.49883, -21.38749, -20.19584, -19.37302, 
    -15.60286, -13.21966, -10.27934, -6.47839, -2.423233, 0.8416929, 
    2.629317, 2.682973, 1.127324, -1.526515, -4.934866, 2.727127, 1.731334, 
    1.399889,
  -33.02792, -32.97892, -32.56007, -31.72274, -30.74157, -30.04212, 
    -26.56238, -22.44532, -16.93535, -10.63038, -5.426571, -2.887532, 
    -3.154822, -5.560196, -9.145553, -12.84596, -16.253, -7.558589, 
    -7.506595, -7.134245,
  -41.52091, -41.82645, -41.99865, -41.91542, -41.78218, -41.88518, 
    -37.62866, -32.77438, -25.59829, -17.70382, -12.13986, -10.84858, 
    -13.45127, -18.29648, -23.40448, -27.10626, -28.9713, -21.69652, 
    -20.11495, -18.93218,
  -46.95891, -47.62904, -48.49966, -49.42086, -50.5189, -51.88708, -46.08807, 
    -41.49573, -34.02331, -25.98105, -21.06019, -21.24872, -25.64825, 
    -31.74947, -36.83765, -39.14276, -38.46293, -34.58241, -31.57569, 
    -29.76226,
  -47.71564, -48.63408, -50.04551, -51.83282, -54.1223, -56.84823, -49.17932, 
    -45.32647, -38.81025, -32.06816, -28.64524, -30.133, -35.16269, 
    -40.78548, -44.25817, -44.35388, -41.14304, -41.3553, -37.41594, -35.31955,
  -43.26765, -44.18139, -45.70936, -47.89296, -51.07134, -55.11771, 
    -45.28218, -41.74169, -36.57541, -31.92972, -30.45863, -32.9719, 
    -37.75286, -41.90597, -43.21301, -41.22623, -36.04288, -39.82709, 
    -35.27989, -33.17536,
  -34.90863, -35.59193, -36.77063, -38.54211, -41.24631, -44.77388, 
    -35.19663, -32.60701, -28.84245, -25.64018, -24.91381, -27.07379, 
    -30.68512, -33.54626, -34.07974, -32.03696, -27.33021, -32.72275, 
    -28.90763, -27.21598,
  -23.41607, -23.71983, -24.23236, -25.01921, -26.24831, -27.88484, 
    -22.12504, -20.9794, -18.80038, -16.65626, -15.81377, -16.65523, 
    -18.51581, -20.25143, -20.92306, -20.17303, -17.7497, -22.14219, 
    -20.23015, -19.32695,
  -9.222198, -9.051055, -8.756757, -8.487967, -8.437077, -8.691723, -7.38933, 
    -7.215876, -6.626178, -5.777412, -5.001366, -4.583436, -4.683494, 
    -5.281631, -6.125695, -6.836977, -7.0343, -8.702703, -8.553235, -8.471096,
  2.890168, 2.81808, 2.673615, 2.529935, 2.493084, 2.578595, 2.801432, 
    2.251043, 1.391916, 0.3291157, -0.7221813, -1.500882, -1.813942, 
    -1.619744, -1.051959, -0.349914, 0.2457331, 0.2097199, 0.2388732, 
    0.1701171,
  5.633145, 6.038826, 6.585892, 7.142332, 7.730578, 8.245561, 8.968597, 
    6.471315, 3.2375, -0.04772019, -2.575249, -3.744222, -3.509316, 
    -2.368634, -1.063603, -0.1796885, 0.000436306, -2.128373, -3.353518, 
    -4.299027,
  6.593079, 7.437188, 8.607376, 9.782068, 10.92312, 11.84556, 13.11227, 
    8.715072, 3.147704, -2.311891, -6.21563, -7.632521, -6.711727, -4.509979, 
    -2.367185, -1.207827, -1.371549, -5.584272, -7.923901, -9.619017,
  5.467204, 6.664538, 8.3173, 9.949989, 11.50571, 12.76529, 14.83601, 
    8.622646, 0.8787537, -6.58207, -11.6562, -13.10647, -11.32732, -7.939667, 
    -4.849131, -3.277623, -3.593103, -10.10366, -13.23079, -15.43041,
  2.718457, 4.133296, 6.058751, 7.929542, 9.725857, 11.19009, 14.84213, 
    6.882899, -2.684271, -11.71083, -17.55494, -18.76648, -16.03079, 
    -11.47311, -7.439894, -5.312268, -5.396101, -15.02254, -18.38118, 
    -20.71944,
  -0.7426267, 0.7095222, 2.650192, 4.530863, 6.445705, 8.015826, 14.94425, 
    5.279279, -5.529923, -15.34156, -21.30845, -21.97333, -18.3397, 
    -12.87292, -8.096805, -5.295572, -4.641665, -19.24957, -22.27896, 
    -24.34553,
  -2.899957, -1.626529, -0.03891325, 1.323487, 2.574806, 3.296831, 14.15716, 
    4.170152, -6.509364, -15.92197, -21.26063, -21.26206, -17.23201, 
    -11.69773, -6.915895, -3.743967, -2.034044, -19.64768, -21.13634, 
    -22.48058,
  -2.731282, -1.791395, -0.7932439, -0.2632165, -0.1459572, -0.7434976, 
    10.9336, 2.650995, -6.201447, -13.84136, -17.69184, -16.86766, -12.93015, 
    -8.219767, -4.370599, -1.609579, 0.6797466, -13.92822, -13.87893, 
    -14.59453,
  -0.9377924, -0.3527196, 0.1226422, 0.06737131, -0.475214, -1.717204, 
    7.378398, 1.201578, -5.20419, -10.2895, -12.01432, -10.01344, -5.993457, 
    -2.029219, 0.7654247, 2.595011, 4.323551, -3.250262, -3.09501, -3.673578,
  1.629534, 1.929811, 2.067144, 1.717359, 0.8384306, -0.7925972, 3.864222, 
    -0.2520339, -4.107887, -6.390203, -5.806819, -2.53889, 1.768305, 
    5.397588, 7.542175, 8.46635, 8.926825, 9.868388, 9.464624, 8.808273,
  3.490702, 3.591268, 3.572377, 3.179994, 2.217885, 0.366586, 0.1041341, 
    -2.118709, -3.511692, -3.043001, -0.3027251, 4.030158, 8.587304, 
    12.10297, 13.91081, 14.06245, 12.96718, 22.09782, 20.95605, 20.18352,
  3.07992, 3.014091, 2.903444, 2.5783, 1.721691, -0.06259346, -4.400949, 
    -4.707374, -3.60326, -0.4897587, 4.082458, 9.010042, 13.34736, 16.36955, 
    17.55716, 16.77123, 14.13748, 29.79915, 28.08007, 27.28681,
  -0.4796867, -0.7382965, -1.012705, -1.341475, -2.037661, -3.452022, 
    -10.0281, -8.283871, -4.623496, 0.9065256, 6.793986, 11.59596, 14.83556, 
    16.41003, 16.16208, 14.10101, 10.4066, 30.03814, 28.30362, 27.74017,
  -6.703052, -7.203838, -7.788765, -8.336419, -9.031157, -10.0361, -16.6056, 
    -12.91344, -6.986189, 0.3541079, 6.764966, 10.57771, 11.75451, 10.88504, 
    8.510214, 5.237806, 1.63269, 22.1217, 21.27178, 21.2798,
  -13.70138, -14.46442, -15.47908, -16.49364, -17.53381, -18.51045, 
    -23.00119, -17.90347, -10.56271, -2.495414, 3.432792, 5.497597, 4.060045, 
    0.4590654, -3.817202, -7.399651, -9.367896, 8.714803, 9.591413, 10.41456,
  -18.98097, -19.94841, -21.37899, -22.99309, -24.76418, -26.3992, -27.20296, 
    -21.43359, -13.8382, -6.338771, -1.842941, -1.881977, -5.705883, 
    -11.25971, -16.20231, -18.76583, -18.01944, -5.015965, -2.016101, 
    -0.3587646,
  -20.5826, -21.58735, -23.22773, -25.38244, -28.18453, -31.20376, -26.79213, 
    -20.62669, -13.50813, -7.493468, -4.985362, -7.023492, -12.48367, 
    -18.82109, -23.26505, -24.15275, -20.66505, -14.14356, -8.925332, 
    -6.536244,
  -18.58064, -19.39539, -20.78774, -22.73203, -25.41147, -28.51807, 
    -21.23217, -16.57204, -11.13295, -6.776063, -5.379655, -7.612461, 
    -12.39739, -17.5252, -20.7218, -20.74978, -16.89118, -16.45036, 
    -11.32508, -9.062169,
  -13.19073, -13.63308, -14.39203, -15.45725, -16.92312, -18.70774, 
    -13.65673, -11.55948, -8.593723, -5.95274, -4.890079, -5.866262, 
    -8.302781, -10.99951, -12.73496, -12.77657, -10.55683, -12.53682, -9.833, 
    -8.589915,
  -4.750134, -4.736323, -4.764349, -4.957309, -5.425515, -6.149175, -5.26367, 
    -5.059452, -4.414222, -3.567738, -2.824295, -2.37032, -2.257102, 
    -2.476457, -2.94505, -3.44083, -3.545211, -4.723301, -4.432084, -4.303707,
  -0.7949679, -0.7290056, -0.6083056, -0.3958577, -0.05297649, 0.3625348, 
    0.8145561, 0.383816, -0.4446023, -1.546948, -2.716424, -3.725163, 
    -4.398774, -4.64779, -4.491026, -4.058528, -3.567768, -3.60633, 
    -3.515617, -3.532481,
  -2.984875, -2.427505, -1.605371, -0.70825, 0.2127521, 1.000114, 1.905358, 
    -0.5558336, -3.893718, -7.410374, -10.27989, -11.88625, -12.14127, 
    -11.44233, -10.41175, -9.583401, -9.311913, -11.36997, -12.43486, 
    -13.26425,
  -5.865497, -4.89, -3.483987, -2.022445, -0.6026769, 0.5559297, 2.113123, 
    -2.24347, -7.911548, -13.66044, -18.04968, -20.1078, -19.87245, 
    -18.21263, -16.29307, -14.99591, -14.80264, -18.92127, -20.92353, 
    -22.40379,
  -9.163703, -7.893562, -6.096825, -4.265342, -2.476885, -0.983274, 1.700274, 
    -4.378547, -12.06118, -19.70308, -25.29616, -27.57269, -26.74331, 
    -24.11396, -21.2976, -19.42719, -19.05806, -25.5787, -28.15663, -30.03827,
  -12.14151, -10.73278, -8.776976, -6.79577, -4.782351, -3.05135, 1.663381, 
    -6.040311, -15.31322, -24.31474, -30.62424, -32.79868, -31.27563, 
    -27.72781, -24.06164, -21.49165, -20.5654, -30.41452, -33.14173, -35.13164,
  -13.99237, -12.61337, -10.72655, -8.777144, -6.619673, -4.733643, 3.47458, 
    -5.867491, -16.2445, -25.88974, -32.2804, -34.00262, -31.75942, 
    -27.44948, -23.03135, -19.57321, -17.61987, -32.40343, -35.09455, 
    -36.96674,
  -13.09759, -11.95386, -10.49666, -9.112898, -7.600042, -6.457311, 5.630576, 
    -3.889865, -14.03588, -23.19756, -28.90211, -29.93781, -27.30612, 
    -22.98307, -18.67606, -15.01738, -12.23065, -29.95144, -31.23345, 
    -32.43307,
  -8.872585, -8.09832, -7.292171, -6.806522, -6.466626, -6.613175, 6.023352, 
    -1.746986, -10.09915, -17.5009, -21.63207, -21.64454, -18.85185, 
    -15.20177, -11.96047, -9.169502, -6.402026, -21.20197, -20.78476, 
    -21.26009,
  -2.293597, -1.882849, -1.63797, -1.830118, -2.317616, -3.351019, 5.821678, 
    -0.1716177, -6.392092, -11.42237, -13.40476, -12.00145, -8.7356, 
    -5.436327, -3.02245, -1.181415, 0.8684886, -6.546676, -5.950524, -6.276498,
  5.578632, 5.692926, 5.527452, 4.854658, 3.706015, 1.839344, 5.273725, 
    0.8223199, -3.267244, -5.72695, -5.387036, -2.451534, 1.542037, 4.995646, 
    7.171038, 8.367846, 9.310635, 11.31711, 11.37455, 10.93734,
  13.02796, 12.92652, 12.50817, 11.5485, 9.90838, 7.298741, 4.27087, 
    1.195322, -0.8176872, -0.7318064, 1.799095, 6.086169, 10.79357, 14.66922, 
    17.0219, 17.85188, 17.51427, 29.12791, 28.35176, 27.70041,
  18.06794, 17.80082, 17.23276, 16.15854, 14.29921, 11.34131, 2.63027, 
    1.111828, 1.309789, 3.878688, 8.290588, 13.47309, 18.46008, 22.45141, 
    24.79171, 25.12409, 23.39344, 43.27967, 41.59973, 40.72245,
  19.12691, 18.70702, 18.02304, 16.95776, 15.20665, 12.52609, 0.1343646, 
    0.6018224, 3.221787, 8.107946, 13.90668, 19.27797, 23.7001, 26.90467, 
    28.41702, 27.74803, 24.70043, 50.35152, 48.04607, 47.08649,
  15.82362, 15.24313, 14.41791, 13.38712, 11.94574, 10.03085, -3.347744, 
    -0.5947804, 4.40055, 11.13398, 17.58827, 22.2733, 25.08544, 26.32837, 
    25.98087, 23.87186, 20.11293, 48.20218, 46.07951, 45.38829,
  9.369065, 8.621003, 7.592027, 6.485933, 5.245653, 4.044686, -7.517156, 
    -2.640999, 4.195691, 11.9163, 18.10333, 21.23518, 21.54218, 19.92136, 
    17.12686, 13.76608, 10.58592, 37.34454, 36.62242, 36.65733,
  2.189144, 1.296411, 0.01455688, -1.374802, -2.85824, -4.061235, -11.27055, 
    -4.88791, 2.867252, 10.48554, 15.49337, 16.48329, 13.94949, 9.388686, 
    4.520112, 0.856246, -0.2917299, 21.48279, 23.3174, 24.44061,
  -3.124312, -4.074872, -5.579389, -7.463519, -9.803929, -12.07064, 
    -12.41104, -5.075687, 2.827206, 9.465117, 12.69995, 11.44237, 6.4281, 
    -0.3412495, -6.326417, -9.39972, -7.891805, 6.050996, 11.23733, 13.64083,
  -5.703659, -6.511373, -7.855319, -9.649977, -12.02694, -14.6322, -9.90867, 
    -4.215977, 2.031923, 7.03093, 9.012211, 7.183271, 2.296216, -3.760732, 
    -8.654139, -10.55381, -8.002439, -3.069259, 2.720335, 5.308744,
  -5.084531, -5.569548, -6.382856, -7.468287, -8.904823, -10.62492, 
    -6.543443, -3.927962, -0.5401826, 2.412389, 3.71501, 2.843411, 0.2489848, 
    -2.956957, -5.472474, -6.295083, -4.517465, -4.504337, -1.324685, 
    0.1328797,
  -1.306764, -1.422848, -1.686074, -2.161645, -2.888842, -3.804895, 
    -3.227554, -2.972517, -2.278323, -1.421556, -0.6997379, -0.271898, 
    -0.1338536, -0.2267089, -0.4887809, -0.7943686, -0.7745719, -1.455512, 
    -1.055968, -0.8982434,
  -4.348464, -4.144964, -3.77705, -3.263221, -2.632801, -1.990937, -1.372645, 
    -1.715749, -2.493126, -3.575378, -4.770998, -5.889002, -6.792717, 
    -7.388072, -7.617749, -7.493149, -7.154756, -7.239266, -7.08037, -7.034297,
  -11.15159, -10.50818, -9.539022, -8.473406, -7.396727, -6.4739, -5.384732, 
    -7.779902, -11.09448, -14.66475, -17.69067, -19.57226, -20.2038, 
    -19.89599, -19.13577, -18.35169, -17.91217, -19.8683, -20.6573, -21.30547,
  -17.41201, -16.41146, -14.96197, -13.44696, -11.96023, -10.70783, -8.80777, 
    -13.04443, -18.59946, -24.34683, -28.91395, -31.34903, -31.63282, 
    -30.47076, -28.81499, -27.40891, -26.78231, -30.78315, -32.31225, 
    -33.50486,
  -22.38144, -21.14741, -19.39502, -17.58004, -15.74374, -14.14, -10.81346, 
    -16.67335, -24.06247, -31.5307, -37.21349, -39.89622, -39.71428, 
    -37.74075, -35.28082, -33.2513, -32.24833, -38.79587, -40.78301, -42.32172,
  -25.25782, -23.92561, -22.055, -20.08961, -17.97453, -16.0736, -10.42272, 
    -17.82937, -26.64558, -35.28653, -41.55843, -44.12035, -43.3311, 
    -40.57608, -37.36356, -34.60819, -32.90596, -42.94455, -45.17724, 
    -46.88216,
  -25.51712, -24.21478, -22.38231, -20.36875, -18.00943, -15.88351, 
    -6.793406, -15.80998, -25.69746, -34.91563, -41.21716, -43.32707, 
    -41.86438, -38.39995, -34.42678, -30.66429, -27.78648, -42.48395, 
    -45.12353, -46.96055,
  -21.99024, -20.91212, -19.46846, -17.93687, -16.10209, -14.57182, -1.87365, 
    -11.00083, -20.66227, -29.41199, -35.04406, -36.48169, -34.62827, 
    -31.15018, -27.34159, -23.53282, -20.09093, -37.53718, -38.99272, 
    -40.25217,
  -14.45229, -13.73342, -12.91803, -12.24272, -11.50699, -11.15386, 1.849977, 
    -5.541506, -13.49405, -20.59375, -24.73356, -25.1539, -23.04933, 
    -20.13297, -17.42569, -14.7995, -11.89794, -26.60869, -26.21614, -26.6399,
  -4.033418, -3.670569, -3.418954, -3.450619, -3.607436, -4.238465, 4.730961, 
    -1.087586, -7.150448, -12.11549, -14.27602, -13.32442, -10.64257, 
    -7.878528, -5.825331, -4.103456, -1.974249, -9.167368, -8.410501, 
    -8.610518,
  8.1231, 8.166135, 7.931097, 7.271444, 6.246578, 4.552039, 6.944951, 2.3927, 
    -1.81649, -4.467356, -4.479568, -2.032851, 1.479343, 4.597703, 6.649861, 
    7.955825, 9.214207, 12.04801, 12.46559, 12.21624,
  20.23377, 20.01342, 19.39205, 18.20719, 16.378, 13.61926, 8.479969, 
    5.021244, 2.63516, 2.315351, 4.378143, 8.199257, 12.56373, 16.31936, 
    18.82285, 20.07989, 20.41599, 33.93286, 33.65987, 33.22082,
  30.12721, 29.70125, 28.80643, 27.26981, 24.89258, 21.43346, 9.357199, 
    7.205256, 6.811886, 8.813684, 12.72072, 17.55532, 22.43349, 26.61425, 
    29.47231, 30.60849, 29.86487, 53.09265, 51.87957, 51.14301,
  35.80163, 35.22631, 34.18043, 32.53546, 30.05577, 26.6112, 9.530968, 
    9.208608, 11.07284, 15.29064, 20.63651, 25.89499, 30.58678, 34.45009, 
    36.97006, 37.46573, 35.4594, 66.05766, 63.86562, 62.82766,
  36.15244, 35.47931, 34.39089, 32.86997, 30.73586, 28.04219, 8.805143, 
    10.81259, 15.01411, 21.08367, 27.24429, 32.16191, 35.73864, 38.20187, 
    39.33059, 38.50361, 35.33881, 69.90232, 67.22041, 66.12025,
  31.5382, 30.80077, 29.71376, 28.39981, 26.77437, 25.10784, 6.990651, 
    11.45378, 17.68668, 24.92493, 31.09442, 34.84584, 36.36159, 36.32405, 
    35.06025, 32.51173, 28.92345, 63.33121, 61.38042, 60.7428,
  23.81192, 23.02013, 21.88388, 20.6134, 19.17506, 18.0226, 4.3634, 10.88234, 
    18.473, 25.99112, 31.33699, 33.23861, 32.0409, 28.83737, 24.75102, 
    20.7322, 18.01102, 47.86461, 48.36767, 48.85758,
  15.65544, 14.81453, 13.51164, 11.9045, 9.922823, 8.159437, 2.46928, 
    10.41016, 18.6689, 25.6863, 29.60525, 29.35598, 25.38231, 19.12127, 
    12.54126, 7.683562, 6.816936, 27.95453, 32.61668, 34.84539,
  8.668119, 7.928811, 6.727989, 5.160435, 3.103199, 0.9296985, 2.266694, 
    8.582815, 15.3137, 20.79737, 23.42366, 22.33655, 17.98784, 11.8105, 
    5.832978, 2.109327, 2.813999, 12.41731, 18.47009, 21.2465,
  4.114567, 3.626065, 2.826355, 1.79008, 0.4242077, -1.222187, 1.360662, 
    4.302523, 7.955643, 11.16317, 12.78221, 12.23697, 9.822134, 6.459996, 
    3.379914, 1.748438, 2.835122, 5.102051, 8.588825, 10.19531,
  2.490541, 2.234663, 1.740663, 1.020608, 0.09634221, -0.9531718, -0.7759612, 
    -0.4986989, 0.2162496, 1.081035, 1.808321, 2.244152, 2.410998, 2.405059, 
    2.309735, 2.207268, 2.399994, 2.389263, 2.914076, 3.103595,
  -7.460973, -7.135199, -6.561992, -5.820375, -4.990794, -4.196261, 
    -3.432629, -3.67939, -4.358079, -5.346859, -6.474012, -7.583599, 
    -8.58357, -9.40663, -9.968849, -10.18909, -10.09926, -10.34927, 
    -10.18853, -10.10984,
  -18.17853, -17.51646, -16.519, -15.42167, -14.30046, -13.29776, -11.95471, 
    -14.19566, -17.32288, -20.73866, -23.69624, -25.63916, -26.47896, 
    -26.47828, -26.00764, -25.35948, -24.84066, -26.8197, -27.35113, -27.82395,
  -27.15875, -26.21721, -24.86359, -23.44147, -21.99411, -20.69617, 
    -18.36661, -22.38428, -27.62712, -33.09493, -37.51141, -39.99078, 
    -40.52509, -39.72727, -38.36655, -36.99676, -36.08423, -40.14152, 
    -41.25758, -42.19146,
  -33.3134, -32.17501, -30.5633, -28.8655, -27.06391, -25.41308, -21.45948, 
    -27.06675, -34.02589, -41.05795, -46.44715, -49.08418, -49.13137, 
    -47.55237, -45.42214, -43.40769, -42.01618, -48.78271, -50.36015, 
    -51.64742,
  -35.92424, -34.67458, -32.90139, -30.97861, -28.82257, -26.84949, 
    -20.49593, -27.66609, -36.00804, -44.10349, -49.95458, -52.37071, 
    -51.75942, -49.3925, -46.51517, -43.74541, -41.59565, -51.90684, 
    -53.95579, -55.53778,
  -34.81084, -33.5298, -31.67455, -29.55705, -27.05094, -24.82203, -15.32626, 
    -24.1346, -33.61255, -42.29888, -48.15695, -50.09172, -48.78105, 
    -45.67623, -41.9831, -38.10069, -34.67702, -49.14528, -52.06219, -54.06459,
  -29.21849, -28.10051, -26.51789, -24.73264, -22.59879, -20.8267, -8.154384, 
    -17.06039, -26.37303, -34.6613, -39.92396, -41.257, -39.59541, -36.48343, 
    -32.97274, -29.14258, -25.38037, -42.24994, -44.23171, -45.76519,
  -19.18343, -18.38516, -17.3571, -16.32338, -15.14655, -14.38697, -1.611324, 
    -8.807798, -16.48705, -23.26277, -27.21244, -27.69538, -25.86983, 
    -23.3253, -20.94514, -18.49685, -15.66615, -29.9958, -30.00192, -30.57594,
  -5.897764, -5.438786, -4.951236, -4.598796, -4.28278, -4.466563, 3.985432, 
    -1.713078, -7.650914, -12.53006, -14.78354, -14.14172, -11.87545, 
    -9.491993, -7.704247, -6.114242, -4.040985, -10.90399, -10.26757, -10.4851,
  9.489427, 9.599062, 9.536472, 9.178855, 8.558449, 7.289674, 8.730269, 
    4.232626, 2.43187e-05, -2.817808, -3.218725, -1.336338, 1.600402, 
    4.28902, 6.1287, 7.444036, 8.890964, 12.36602, 13.00596, 12.8882,
  25.2313, 25.00916, 24.42213, 23.35938, 21.76686, 19.33428, 12.60745, 
    9.130114, 6.582012, 5.879066, 7.325941, 10.40671, 14.08389, 17.36551, 
    19.70704, 21.15604, 22.029, 36.90626, 37.19161, 37.02418,
  39.13785, 38.63342, 37.61174, 35.97002, 33.58445, 30.24705, 15.71522, 
    13.42562, 12.72129, 14.17588, 17.35349, 21.41488, 25.62547, 29.38802, 
    32.2091, 33.7717, 33.91663, 59.5942, 59.16719, 58.77601,
  49.01458, 48.31395, 47.02538, 45.07981, 42.3328, 38.72884, 18.12319, 
    17.50261, 18.89756, 22.46616, 27.10326, 31.73704, 35.98342, 39.68225, 
    42.44649, 43.65531, 42.75574, 77.14975, 75.7072, 74.94414,
  53.27028, 52.48289, 51.1397, 49.2402, 46.66997, 43.57441, 19.68046, 
    21.26591, 24.88529, 30.2962, 35.91215, 40.53904, 44.11454, 46.89465, 
    48.69989, 48.82584, 46.63726, 86.40283, 84.03204, 82.95117,
  51.46915, 50.68752, 49.45321, 47.84952, 45.80912, 43.69381, 19.99628, 
    24.06657, 29.74064, 36.44886, 42.3762, 46.30996, 48.41254, 49.27863, 
    49.0802, 47.41948, 44.10769, 84.90311, 82.50626, 81.53608,
  44.59925, 43.85416, 42.73905, 41.38968, 39.7554, 38.37519, 18.77499, 
    25.12642, 32.37617, 39.65568, 45.16196, 47.74332, 47.65779, 45.73913, 
    42.68142, 38.88176, 35.20739, 72.0328, 71.48416, 71.43936,
  34.8574, 34.10093, 32.91765, 31.41747, 29.53897, 27.9327, 16.77654, 
    24.81431, 33.07148, 40.24849, 44.74447, 45.5481, 42.91704, 37.82816, 
    31.59097, 25.72564, 22.58687, 50.15359, 53.9406, 55.85922,
  24.09682, 23.42819, 22.34345, 20.90891, 19.00482, 17.0389, 14.38952, 
    20.89367, 27.76996, 33.5507, 36.8087, 36.68118, 33.39294, 27.91995, 
    21.75649, 16.72346, 15.36221, 29.5211, 35.31533, 38.08797,
  14.25819, 13.7781, 12.99523, 11.97338, 10.59863, 8.933764, 9.483008, 
    12.51692, 16.23907, 19.60618, 21.58067, 21.56398, 19.70165, 16.67012, 
    13.47446, 11.24934, 11.50743, 16.24285, 19.76069, 21.40061,
  6.561945, 6.169615, 5.462528, 4.529089, 3.434735, 2.264529, 1.909531, 
    2.150112, 2.832741, 3.686478, 4.444645, 4.951902, 5.221179, 5.349418, 
    5.43445, 5.550624, 5.94936, 6.792755, 7.459654, 7.690007,
  -10.70534, -10.24702, -9.465092, -8.508974, -7.497489, -6.550989, 
    -5.575246, -5.652989, -6.111263, -6.844917, -7.708451, -8.593334, 
    -9.479903, -10.37931, -11.25296, -11.97989, -12.45516, -13.29091, 
    -13.42783, -13.47643,
  -25.32955, -24.70602, -23.76875, -22.71719, -21.57674, -20.45534, 
    -18.61446, -20.51123, -23.14337, -26.01205, -28.45841, -30.02456, 
    -30.72065, -30.84731, -30.71325, -30.45237, -30.19728, -32.73788, 
    -33.27361, -33.70723,
  -36.9234, -36.10928, -34.95018, -33.69981, -32.31636, -30.95064, -27.91145, 
    -31.53461, -36.11628, -40.8097, -44.47894, -46.38593, -46.65358, 
    -45.92148, -44.84256, -43.7425, -42.88599, -47.63251, -48.66134, -49.51094,
  -44.11095, -43.09494, -41.65901, -40.10888, -38.37254, -36.72737, 
    -32.01044, -37.31032, -43.58286, -49.70896, -54.15956, -56.02339, 
    -55.62793, -53.97257, -51.99953, -50.11617, -48.63014, -56.19534, 
    -57.82533, -59.11663,
  -46.35525, -45.14574, -43.40794, -41.495, -39.34914, -37.45214, -30.56668, 
    -37.57301, -45.3285, -52.50528, -57.32431, -58.8366, -57.63726, 
    -55.04155, -52.15815, -49.34061, -46.95512, -57.79887, -60.25779, -62.0639,
  -43.88313, -42.50795, -40.47065, -38.16132, -35.58611, -33.47569, 
    -24.16712, -32.88465, -41.95348, -49.84096, -54.72123, -55.75941, 
    -53.82074, -50.39759, -46.5581, -42.44645, -38.63953, -52.53195, 
    -56.31602, -58.8923,
  -36.39621, -35.06542, -33.09743, -30.88808, -28.47235, -26.6429, -14.96738, 
    -23.79346, -32.80375, -40.43188, -44.89274, -45.52686, -43.39721, 
    -40.05171, -36.43253, -32.4528, -28.5237, -43.98286, -47.15054, -49.39227,
  -24.14521, -23.0539, -21.49063, -19.81939, -18.07751, -16.95271, -5.413638, 
    -12.55752, -19.99449, -26.29502, -29.77106, -29.9593, -28.02144, 
    -25.47224, -23.12954, -20.7405, -18.11472, -31.21965, -32.31823, -33.4302,
  -8.295929, -7.496875, -6.3853, -5.260063, -4.186494, -3.765842, 3.397103, 
    -2.209377, -7.99539, -12.70102, -14.95646, -14.55665, -12.64309, 
    -10.55938, -8.947614, -7.447442, -5.530171, -11.55362, -11.525, -12.01637,
  10.06204, 10.49782, 11.04704, 11.49388, 11.75026, 11.31556, 11.35391, 
    7.077068, 2.92949, -0.04402536, -0.9569264, 0.1200773, 2.192249, 
    4.195764, 5.650996, 6.881093, 8.441914, 12.66889, 13.34056, 13.27206,
  29.32716, 29.35391, 29.25722, 28.90495, 28.1957, 26.75104, 18.28952, 
    15.16978, 12.64272, 11.48395, 11.98702, 13.8039, 16.17806, 18.39733, 
    20.11804, 21.49549, 22.85878, 38.86724, 39.87074, 40.1013,
  47.44909, 47.0732, 46.33697, 45.19168, 43.54229, 41.16434, 24.2387, 
    22.33496, 21.53741, 22.29163, 24.25458, 26.8116, 29.48653, 31.95573, 
    34.0056, 35.56355, 36.61091, 64.30976, 65.24428, 65.56868,
  62.24054, 61.53976, 60.30015, 58.55505, 56.24039, 53.32462, 29.30364, 
    28.9253, 30.04421, 32.75001, 36.11681, 39.30153, 42.09992, 44.56694, 
    46.62938, 48.00548, 48.35852, 86.12791, 86.4759, 86.60828,
  71.80052, 70.91587, 69.42068, 67.41796, 64.88706, 62.02287, 33.41351, 
    34.97066, 38.11294, 42.6215, 47.15256, 50.71114, 53.31258, 55.32219, 
    56.8115, 57.37508, 56.53413, 101.3328, 100.7001, 100.4232,
  74.88444, 73.97131, 72.48312, 70.56344, 68.22305, 65.8914, 36.14684, 
    39.92439, 44.99551, 50.92296, 56.1809, 59.72202, 61.69623, 62.66193, 
    62.83226, 61.84132, 59.40931, 106.8564, 105.4545, 104.8739,
  71.18228, 70.33372, 68.98109, 67.26654, 65.20522, 63.41928, 36.8078, 
    42.73167, 49.40566, 56.19684, 61.61981, 64.66382, 65.51012, 64.77205, 
    62.81319, 59.57185, 55.48896, 99.9812, 99.18762, 98.98291,
  61.50531, 60.67846, 59.32269, 57.55483, 55.408, 53.5967, 35.15945, 
    42.70986, 50.54302, 57.63936, 62.68756, 64.77808, 64.02946, 60.98133, 
    56.16194, 50.12245, 44.63254, 79.62478, 82.20426, 83.74281,
  47.05713, 46.33891, 45.12409, 43.47293, 41.34857, 39.25682, 30.35932, 
    36.49104, 43.07636, 48.95496, 52.95988, 54.28512, 52.96988, 49.48023, 
    44.47703, 38.9083, 34.97865, 55.28802, 59.95537, 62.44661,
  30.03084, 29.48631, 28.55681, 27.28878, 25.59663, 23.66111, 20.47712, 
    23.27327, 26.76046, 30.1482, 32.59478, 33.5291, 32.94987, 31.19156, 
    28.78527, 26.45987, 25.63287, 34.3974, 37.44922, 38.92793,
  12.70131, 12.13377, 11.1471, 9.91159, 8.542149, 7.157581, 5.786036, 
    5.863673, 6.392272, 7.169528, 7.97947, 8.674801, 9.244339, 9.74291, 
    10.23248, 10.75917, 11.50989, 13.93886, 14.87192, 15.22682,
  -11.63917, -11.13408, -10.28048, -9.251871, -8.176452, -7.171406, 
    -6.079078, -6.062316, -6.372009, -6.906917, -7.531162, -8.161996, 
    -8.826924, -9.599981, -10.50843, -11.47044, -12.35414, -13.75531, 
    -14.32323, -14.6181,
  -27.30098, -26.69423, -25.77779, -24.73112, -23.55918, -22.36731, 
    -20.20902, -21.90314, -24.18815, -26.60343, -28.53317, -29.59085, 
    -29.8835, -29.79776, -29.68661, -29.66043, -29.76277, -33.01524, 
    -33.92859, -34.57604,
  -39.59485, -38.81941, -37.71314, -36.49979, -35.11585, -33.72102, 
    -30.28043, -33.7028, -37.85763, -41.95243, -44.92163, -46.13285, 
    -45.8378, -44.77443, -43.62656, -42.66612, -42.05398, -47.58787, 
    -49.00456, -50.07993,
  -47.06993, -46.07312, -44.66198, -43.13652, -41.43008, -39.84213, 
    -34.80252, -39.99238, -45.8738, -51.36826, -55.03869, -56.10285, 
    -55.02918, -52.91546, -50.72747, -48.81524, -47.41084, -55.65848, 
    -57.74934, -59.31717,
  -49.23507, -47.99784, -46.21674, -44.28439, -42.19109, -40.43953, 
    -33.50888, -40.49791, -47.95993, -54.5539, -58.60321, -59.29942, 
    -57.37199, -54.22306, -50.98096, -47.95529, -45.4897, -56.59233, 
    -59.62409, -61.79155,
  -46.42253, -44.95454, -42.77914, -40.38209, -37.86482, -35.95444, -27.1461, 
    -35.85394, -44.73259, -52.13935, -56.33641, -56.62336, -53.97884, 
    -49.96817, -45.6842, -41.25597, -37.2866, -50.55977, -54.97514, -58.01217,
  -38.49254, -37.00623, -34.79332, -32.37263, -29.8949, -28.15631, -17.57704, 
    -26.39145, -35.26555, -42.5026, -46.41536, -46.46464, -43.78083, 
    -39.94917, -35.93767, -31.68444, -27.68591, -41.80426, -45.76243, -48.5232,
  -25.72577, -24.42321, -22.50743, -20.46733, -18.45499, -17.19966, 
    -6.907176, -14.06424, -21.38556, -27.39231, -30.52494, -30.41173, 
    -28.21134, -25.41377, -22.84688, -20.31683, -17.77381, -29.55761, 
    -31.49784, -33.06738,
  -9.210961, -8.148962, -6.587311, -4.952544, -3.425573, -2.66805, 3.3733, 
    -2.192581, -7.881507, -12.44701, -14.63726, -14.28679, -12.46608, 
    -10.43244, -8.8019, -7.26563, -5.432866, -10.57791, -11.11955, -11.90135,
  10.01556, 10.74555, 11.81022, 12.87803, 13.75543, 13.87966, 12.95419, 
    8.848155, 4.799569, 1.794064, 0.6435242, 1.300597, 2.894164, 4.497474, 
    5.70972, 6.854819, 8.407971, 13.09673, 13.59089, 13.44719,
  30.45658, 30.776, 31.20541, 31.52676, 31.55868, 30.87201, 21.51591, 
    18.72273, 16.30089, 14.94256, 14.93056, 16, 17.54465, 19.01884, 20.21659, 
    21.37964, 22.85435, 39.11512, 40.38075, 40.77939,
  50.18473, 50.06216, 49.79597, 49.29362, 48.41444, 46.9, 28.98488, 27.50993, 
    26.79262, 27.19688, 28.43781, 30.02628, 31.63116, 33.09507, 34.39137, 
    35.63259, 36.93675, 64.96223, 66.62106, 67.37151,
  67.10821, 66.58578, 65.69347, 64.46476, 62.8237, 60.71905, 35.40749, 
    35.44323, 36.56585, 38.80814, 41.35868, 43.51492, 45.18253, 46.55063, 
    47.75425, 48.77902, 49.53716, 88.01234, 89.51743, 90.30977,
  79.30547, 78.4995, 77.17686, 75.47682, 73.39426, 71.11259, 40.71096, 
    42.53741, 45.56898, 49.56606, 53.33112, 55.99737, 57.637, 58.69095, 
    59.41317, 59.68872, 59.34621, 105.5035, 106.3032, 106.8156,
  85.26352, 84.32523, 82.81702, 80.94095, 78.746, 76.65497, 44.48794, 
    48.29914, 53.14144, 58.59456, 63.28709, 66.27293, 67.707, 68.14821, 
    67.89941, 66.79022, 64.78082, 114.3846, 114.3314, 114.4658,
  84.04198, 83.08468, 81.54977, 79.64882, 77.46265, 75.61214, 45.95056, 
    51.6445, 57.99641, 64.42953, 69.60615, 72.59215, 73.54076, 72.98575, 
    71.20938, 68.08212, 64.02373, 111.3482, 111.3001, 111.5033,
  75.49812, 74.51241, 72.88265, 70.81219, 68.43785, 66.47202, 44.39825, 
    51.44211, 58.87345, 65.76664, 70.93062, 73.51214, 73.58983, 71.54795, 
    67.60579, 61.85013, 55.60539, 93.74643, 96.02483, 97.57922,
  60.00261, 59.11932, 57.60606, 55.5959, 53.16988, 50.8976, 38.30669, 
    43.96084, 50.16017, 55.91314, 60.18506, 62.22158, 62.01585, 59.84041, 
    55.95539, 50.72466, 45.8033, 69.51892, 73.38236, 75.68821,
  39.34684, 38.67354, 37.49446, 35.88765, 33.84902, 31.67924, 25.96256, 
    28.4901, 31.69341, 34.96492, 37.59253, 39.05034, 39.30038, 38.52928, 
    36.99052, 35.0491, 33.78917, 45.33301, 47.96998, 49.33248,
  16.19508, 15.54678, 14.4164, 13.00132, 11.45139, 9.931472, 7.847852, 
    7.797616, 8.188686, 8.878651, 9.690671, 10.4915, 11.26515, 12.04185, 
    12.84472, 13.67657, 14.66263, 18.25719, 19.44049, 19.97217 ;

 b =
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -30, -30, -30, -30, -30, -30, -30, -30, -30, 
    -30, -30, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50,
  -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, -50, 
    -50, -50, -50, -50, -50 ;
}
